//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][18]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul  7 02:19:44 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__18_ -----
module sb_1__18_(prog_clk,
                 chanx_right_in,
                 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                 right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                 right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                 chany_bottom_in,
                 bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                 bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                 bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                 chanx_left_in,
                 left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                 left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                 left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                 ccff_head,
                 chanx_right_out,
                 chany_bottom_out,
                 chanx_left_out,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:284] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:284] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:284] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:284] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:284] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:284] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_100_sram;
wire [0:2] mux_tree_tapbuf_size4_100_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_101_sram;
wire [0:2] mux_tree_tapbuf_size4_101_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_102_sram;
wire [0:2] mux_tree_tapbuf_size4_102_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_103_sram;
wire [0:2] mux_tree_tapbuf_size4_103_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_104_sram;
wire [0:2] mux_tree_tapbuf_size4_104_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_105_sram;
wire [0:2] mux_tree_tapbuf_size4_105_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_106_sram;
wire [0:2] mux_tree_tapbuf_size4_106_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_107_sram;
wire [0:2] mux_tree_tapbuf_size4_107_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_108_sram;
wire [0:2] mux_tree_tapbuf_size4_108_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_109_sram;
wire [0:2] mux_tree_tapbuf_size4_109_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_10_sram;
wire [0:2] mux_tree_tapbuf_size4_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_110_sram;
wire [0:2] mux_tree_tapbuf_size4_110_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_111_sram;
wire [0:2] mux_tree_tapbuf_size4_111_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_112_sram;
wire [0:2] mux_tree_tapbuf_size4_112_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_113_sram;
wire [0:2] mux_tree_tapbuf_size4_113_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_114_sram;
wire [0:2] mux_tree_tapbuf_size4_114_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_115_sram;
wire [0:2] mux_tree_tapbuf_size4_115_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_116_sram;
wire [0:2] mux_tree_tapbuf_size4_116_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_117_sram;
wire [0:2] mux_tree_tapbuf_size4_117_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_118_sram;
wire [0:2] mux_tree_tapbuf_size4_118_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_119_sram;
wire [0:2] mux_tree_tapbuf_size4_119_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_11_sram;
wire [0:2] mux_tree_tapbuf_size4_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_120_sram;
wire [0:2] mux_tree_tapbuf_size4_120_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_121_sram;
wire [0:2] mux_tree_tapbuf_size4_121_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_122_sram;
wire [0:2] mux_tree_tapbuf_size4_122_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_123_sram;
wire [0:2] mux_tree_tapbuf_size4_123_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_124_sram;
wire [0:2] mux_tree_tapbuf_size4_124_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_125_sram;
wire [0:2] mux_tree_tapbuf_size4_125_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_126_sram;
wire [0:2] mux_tree_tapbuf_size4_126_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_127_sram;
wire [0:2] mux_tree_tapbuf_size4_127_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_128_sram;
wire [0:2] mux_tree_tapbuf_size4_128_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_129_sram;
wire [0:2] mux_tree_tapbuf_size4_129_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_12_sram;
wire [0:2] mux_tree_tapbuf_size4_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_130_sram;
wire [0:2] mux_tree_tapbuf_size4_130_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_131_sram;
wire [0:2] mux_tree_tapbuf_size4_131_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_132_sram;
wire [0:2] mux_tree_tapbuf_size4_132_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_133_sram;
wire [0:2] mux_tree_tapbuf_size4_133_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_134_sram;
wire [0:2] mux_tree_tapbuf_size4_134_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_135_sram;
wire [0:2] mux_tree_tapbuf_size4_135_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_136_sram;
wire [0:2] mux_tree_tapbuf_size4_136_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_137_sram;
wire [0:2] mux_tree_tapbuf_size4_137_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_138_sram;
wire [0:2] mux_tree_tapbuf_size4_138_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_139_sram;
wire [0:2] mux_tree_tapbuf_size4_139_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_13_sram;
wire [0:2] mux_tree_tapbuf_size4_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_140_sram;
wire [0:2] mux_tree_tapbuf_size4_140_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_141_sram;
wire [0:2] mux_tree_tapbuf_size4_141_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_142_sram;
wire [0:2] mux_tree_tapbuf_size4_142_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_143_sram;
wire [0:2] mux_tree_tapbuf_size4_143_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_144_sram;
wire [0:2] mux_tree_tapbuf_size4_144_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_145_sram;
wire [0:2] mux_tree_tapbuf_size4_145_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_146_sram;
wire [0:2] mux_tree_tapbuf_size4_146_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_147_sram;
wire [0:2] mux_tree_tapbuf_size4_147_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_148_sram;
wire [0:2] mux_tree_tapbuf_size4_148_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_149_sram;
wire [0:2] mux_tree_tapbuf_size4_149_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_14_sram;
wire [0:2] mux_tree_tapbuf_size4_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_150_sram;
wire [0:2] mux_tree_tapbuf_size4_150_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_151_sram;
wire [0:2] mux_tree_tapbuf_size4_151_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_152_sram;
wire [0:2] mux_tree_tapbuf_size4_152_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_153_sram;
wire [0:2] mux_tree_tapbuf_size4_153_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_154_sram;
wire [0:2] mux_tree_tapbuf_size4_154_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_155_sram;
wire [0:2] mux_tree_tapbuf_size4_155_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_156_sram;
wire [0:2] mux_tree_tapbuf_size4_156_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_157_sram;
wire [0:2] mux_tree_tapbuf_size4_157_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_158_sram;
wire [0:2] mux_tree_tapbuf_size4_158_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_159_sram;
wire [0:2] mux_tree_tapbuf_size4_159_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_15_sram;
wire [0:2] mux_tree_tapbuf_size4_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_160_sram;
wire [0:2] mux_tree_tapbuf_size4_160_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_161_sram;
wire [0:2] mux_tree_tapbuf_size4_161_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_162_sram;
wire [0:2] mux_tree_tapbuf_size4_162_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_163_sram;
wire [0:2] mux_tree_tapbuf_size4_163_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_164_sram;
wire [0:2] mux_tree_tapbuf_size4_164_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_165_sram;
wire [0:2] mux_tree_tapbuf_size4_165_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_166_sram;
wire [0:2] mux_tree_tapbuf_size4_166_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_167_sram;
wire [0:2] mux_tree_tapbuf_size4_167_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_168_sram;
wire [0:2] mux_tree_tapbuf_size4_168_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_169_sram;
wire [0:2] mux_tree_tapbuf_size4_169_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_16_sram;
wire [0:2] mux_tree_tapbuf_size4_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_170_sram;
wire [0:2] mux_tree_tapbuf_size4_170_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_171_sram;
wire [0:2] mux_tree_tapbuf_size4_171_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_172_sram;
wire [0:2] mux_tree_tapbuf_size4_172_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_173_sram;
wire [0:2] mux_tree_tapbuf_size4_173_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_174_sram;
wire [0:2] mux_tree_tapbuf_size4_174_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_175_sram;
wire [0:2] mux_tree_tapbuf_size4_175_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_176_sram;
wire [0:2] mux_tree_tapbuf_size4_176_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_177_sram;
wire [0:2] mux_tree_tapbuf_size4_177_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_178_sram;
wire [0:2] mux_tree_tapbuf_size4_178_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_179_sram;
wire [0:2] mux_tree_tapbuf_size4_179_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_17_sram;
wire [0:2] mux_tree_tapbuf_size4_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_180_sram;
wire [0:2] mux_tree_tapbuf_size4_180_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_181_sram;
wire [0:2] mux_tree_tapbuf_size4_181_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_182_sram;
wire [0:2] mux_tree_tapbuf_size4_182_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_183_sram;
wire [0:2] mux_tree_tapbuf_size4_183_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_184_sram;
wire [0:2] mux_tree_tapbuf_size4_184_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_185_sram;
wire [0:2] mux_tree_tapbuf_size4_185_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_186_sram;
wire [0:2] mux_tree_tapbuf_size4_186_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_187_sram;
wire [0:2] mux_tree_tapbuf_size4_187_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_188_sram;
wire [0:2] mux_tree_tapbuf_size4_188_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_189_sram;
wire [0:2] mux_tree_tapbuf_size4_189_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_18_sram;
wire [0:2] mux_tree_tapbuf_size4_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_190_sram;
wire [0:2] mux_tree_tapbuf_size4_190_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_191_sram;
wire [0:2] mux_tree_tapbuf_size4_191_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_192_sram;
wire [0:2] mux_tree_tapbuf_size4_192_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_193_sram;
wire [0:2] mux_tree_tapbuf_size4_193_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_194_sram;
wire [0:2] mux_tree_tapbuf_size4_194_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_195_sram;
wire [0:2] mux_tree_tapbuf_size4_195_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_196_sram;
wire [0:2] mux_tree_tapbuf_size4_196_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_197_sram;
wire [0:2] mux_tree_tapbuf_size4_197_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_198_sram;
wire [0:2] mux_tree_tapbuf_size4_198_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_199_sram;
wire [0:2] mux_tree_tapbuf_size4_199_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_19_sram;
wire [0:2] mux_tree_tapbuf_size4_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_200_sram;
wire [0:2] mux_tree_tapbuf_size4_200_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_201_sram;
wire [0:2] mux_tree_tapbuf_size4_201_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_202_sram;
wire [0:2] mux_tree_tapbuf_size4_202_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_203_sram;
wire [0:2] mux_tree_tapbuf_size4_203_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_204_sram;
wire [0:2] mux_tree_tapbuf_size4_204_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_205_sram;
wire [0:2] mux_tree_tapbuf_size4_205_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_206_sram;
wire [0:2] mux_tree_tapbuf_size4_206_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_207_sram;
wire [0:2] mux_tree_tapbuf_size4_207_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_208_sram;
wire [0:2] mux_tree_tapbuf_size4_208_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_209_sram;
wire [0:2] mux_tree_tapbuf_size4_209_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_20_sram;
wire [0:2] mux_tree_tapbuf_size4_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_210_sram;
wire [0:2] mux_tree_tapbuf_size4_210_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_211_sram;
wire [0:2] mux_tree_tapbuf_size4_211_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_212_sram;
wire [0:2] mux_tree_tapbuf_size4_212_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_213_sram;
wire [0:2] mux_tree_tapbuf_size4_213_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_214_sram;
wire [0:2] mux_tree_tapbuf_size4_214_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_215_sram;
wire [0:2] mux_tree_tapbuf_size4_215_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_216_sram;
wire [0:2] mux_tree_tapbuf_size4_216_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_217_sram;
wire [0:2] mux_tree_tapbuf_size4_217_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_218_sram;
wire [0:2] mux_tree_tapbuf_size4_218_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_219_sram;
wire [0:2] mux_tree_tapbuf_size4_219_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_21_sram;
wire [0:2] mux_tree_tapbuf_size4_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_220_sram;
wire [0:2] mux_tree_tapbuf_size4_220_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_221_sram;
wire [0:2] mux_tree_tapbuf_size4_221_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_222_sram;
wire [0:2] mux_tree_tapbuf_size4_222_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_223_sram;
wire [0:2] mux_tree_tapbuf_size4_223_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_224_sram;
wire [0:2] mux_tree_tapbuf_size4_224_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_225_sram;
wire [0:2] mux_tree_tapbuf_size4_225_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_22_sram;
wire [0:2] mux_tree_tapbuf_size4_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_23_sram;
wire [0:2] mux_tree_tapbuf_size4_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_24_sram;
wire [0:2] mux_tree_tapbuf_size4_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_25_sram;
wire [0:2] mux_tree_tapbuf_size4_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_26_sram;
wire [0:2] mux_tree_tapbuf_size4_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_27_sram;
wire [0:2] mux_tree_tapbuf_size4_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_28_sram;
wire [0:2] mux_tree_tapbuf_size4_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_29_sram;
wire [0:2] mux_tree_tapbuf_size4_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_30_sram;
wire [0:2] mux_tree_tapbuf_size4_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_31_sram;
wire [0:2] mux_tree_tapbuf_size4_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_32_sram;
wire [0:2] mux_tree_tapbuf_size4_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_33_sram;
wire [0:2] mux_tree_tapbuf_size4_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_34_sram;
wire [0:2] mux_tree_tapbuf_size4_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_35_sram;
wire [0:2] mux_tree_tapbuf_size4_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_36_sram;
wire [0:2] mux_tree_tapbuf_size4_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_37_sram;
wire [0:2] mux_tree_tapbuf_size4_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_38_sram;
wire [0:2] mux_tree_tapbuf_size4_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_39_sram;
wire [0:2] mux_tree_tapbuf_size4_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_40_sram;
wire [0:2] mux_tree_tapbuf_size4_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_41_sram;
wire [0:2] mux_tree_tapbuf_size4_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_42_sram;
wire [0:2] mux_tree_tapbuf_size4_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_43_sram;
wire [0:2] mux_tree_tapbuf_size4_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_44_sram;
wire [0:2] mux_tree_tapbuf_size4_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_45_sram;
wire [0:2] mux_tree_tapbuf_size4_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_46_sram;
wire [0:2] mux_tree_tapbuf_size4_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_47_sram;
wire [0:2] mux_tree_tapbuf_size4_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_48_sram;
wire [0:2] mux_tree_tapbuf_size4_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_49_sram;
wire [0:2] mux_tree_tapbuf_size4_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_50_sram;
wire [0:2] mux_tree_tapbuf_size4_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_51_sram;
wire [0:2] mux_tree_tapbuf_size4_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_52_sram;
wire [0:2] mux_tree_tapbuf_size4_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_53_sram;
wire [0:2] mux_tree_tapbuf_size4_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_54_sram;
wire [0:2] mux_tree_tapbuf_size4_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_55_sram;
wire [0:2] mux_tree_tapbuf_size4_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_56_sram;
wire [0:2] mux_tree_tapbuf_size4_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_57_sram;
wire [0:2] mux_tree_tapbuf_size4_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_58_sram;
wire [0:2] mux_tree_tapbuf_size4_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_59_sram;
wire [0:2] mux_tree_tapbuf_size4_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_60_sram;
wire [0:2] mux_tree_tapbuf_size4_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_61_sram;
wire [0:2] mux_tree_tapbuf_size4_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_62_sram;
wire [0:2] mux_tree_tapbuf_size4_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_63_sram;
wire [0:2] mux_tree_tapbuf_size4_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_64_sram;
wire [0:2] mux_tree_tapbuf_size4_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_65_sram;
wire [0:2] mux_tree_tapbuf_size4_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_66_sram;
wire [0:2] mux_tree_tapbuf_size4_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_67_sram;
wire [0:2] mux_tree_tapbuf_size4_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_68_sram;
wire [0:2] mux_tree_tapbuf_size4_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_69_sram;
wire [0:2] mux_tree_tapbuf_size4_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_70_sram;
wire [0:2] mux_tree_tapbuf_size4_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_71_sram;
wire [0:2] mux_tree_tapbuf_size4_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_72_sram;
wire [0:2] mux_tree_tapbuf_size4_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_73_sram;
wire [0:2] mux_tree_tapbuf_size4_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_74_sram;
wire [0:2] mux_tree_tapbuf_size4_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_75_sram;
wire [0:2] mux_tree_tapbuf_size4_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_76_sram;
wire [0:2] mux_tree_tapbuf_size4_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_77_sram;
wire [0:2] mux_tree_tapbuf_size4_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_78_sram;
wire [0:2] mux_tree_tapbuf_size4_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_79_sram;
wire [0:2] mux_tree_tapbuf_size4_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_7_sram;
wire [0:2] mux_tree_tapbuf_size4_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_80_sram;
wire [0:2] mux_tree_tapbuf_size4_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_81_sram;
wire [0:2] mux_tree_tapbuf_size4_81_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_82_sram;
wire [0:2] mux_tree_tapbuf_size4_82_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_83_sram;
wire [0:2] mux_tree_tapbuf_size4_83_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_84_sram;
wire [0:2] mux_tree_tapbuf_size4_84_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_85_sram;
wire [0:2] mux_tree_tapbuf_size4_85_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_86_sram;
wire [0:2] mux_tree_tapbuf_size4_86_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_87_sram;
wire [0:2] mux_tree_tapbuf_size4_87_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_88_sram;
wire [0:2] mux_tree_tapbuf_size4_88_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_89_sram;
wire [0:2] mux_tree_tapbuf_size4_89_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_8_sram;
wire [0:2] mux_tree_tapbuf_size4_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_90_sram;
wire [0:2] mux_tree_tapbuf_size4_90_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_91_sram;
wire [0:2] mux_tree_tapbuf_size4_91_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_92_sram;
wire [0:2] mux_tree_tapbuf_size4_92_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_93_sram;
wire [0:2] mux_tree_tapbuf_size4_93_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_94_sram;
wire [0:2] mux_tree_tapbuf_size4_94_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_95_sram;
wire [0:2] mux_tree_tapbuf_size4_95_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_96_sram;
wire [0:2] mux_tree_tapbuf_size4_96_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_97_sram;
wire [0:2] mux_tree_tapbuf_size4_97_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_98_sram;
wire [0:2] mux_tree_tapbuf_size4_98_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_99_sram;
wire [0:2] mux_tree_tapbuf_size4_99_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_9_sram;
wire [0:2] mux_tree_tapbuf_size4_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_100_sram;
wire [0:2] mux_tree_tapbuf_size6_100_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_101_sram;
wire [0:2] mux_tree_tapbuf_size6_101_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_102_sram;
wire [0:2] mux_tree_tapbuf_size6_102_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_103_sram;
wire [0:2] mux_tree_tapbuf_size6_103_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_104_sram;
wire [0:2] mux_tree_tapbuf_size6_104_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_105_sram;
wire [0:2] mux_tree_tapbuf_size6_105_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_106_sram;
wire [0:2] mux_tree_tapbuf_size6_106_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_107_sram;
wire [0:2] mux_tree_tapbuf_size6_107_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_108_sram;
wire [0:2] mux_tree_tapbuf_size6_108_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_11_sram;
wire [0:2] mux_tree_tapbuf_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_12_sram;
wire [0:2] mux_tree_tapbuf_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_13_sram;
wire [0:2] mux_tree_tapbuf_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_14_sram;
wire [0:2] mux_tree_tapbuf_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_15_sram;
wire [0:2] mux_tree_tapbuf_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_16_sram;
wire [0:2] mux_tree_tapbuf_size6_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_17_sram;
wire [0:2] mux_tree_tapbuf_size6_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_18_sram;
wire [0:2] mux_tree_tapbuf_size6_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_19_sram;
wire [0:2] mux_tree_tapbuf_size6_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_20_sram;
wire [0:2] mux_tree_tapbuf_size6_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_21_sram;
wire [0:2] mux_tree_tapbuf_size6_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_22_sram;
wire [0:2] mux_tree_tapbuf_size6_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_23_sram;
wire [0:2] mux_tree_tapbuf_size6_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_24_sram;
wire [0:2] mux_tree_tapbuf_size6_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_25_sram;
wire [0:2] mux_tree_tapbuf_size6_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_26_sram;
wire [0:2] mux_tree_tapbuf_size6_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_27_sram;
wire [0:2] mux_tree_tapbuf_size6_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_28_sram;
wire [0:2] mux_tree_tapbuf_size6_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_29_sram;
wire [0:2] mux_tree_tapbuf_size6_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_30_sram;
wire [0:2] mux_tree_tapbuf_size6_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_31_sram;
wire [0:2] mux_tree_tapbuf_size6_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_32_sram;
wire [0:2] mux_tree_tapbuf_size6_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_33_sram;
wire [0:2] mux_tree_tapbuf_size6_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_34_sram;
wire [0:2] mux_tree_tapbuf_size6_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_35_sram;
wire [0:2] mux_tree_tapbuf_size6_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_36_sram;
wire [0:2] mux_tree_tapbuf_size6_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_37_sram;
wire [0:2] mux_tree_tapbuf_size6_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_38_sram;
wire [0:2] mux_tree_tapbuf_size6_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_39_sram;
wire [0:2] mux_tree_tapbuf_size6_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_40_sram;
wire [0:2] mux_tree_tapbuf_size6_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_41_sram;
wire [0:2] mux_tree_tapbuf_size6_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_42_sram;
wire [0:2] mux_tree_tapbuf_size6_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_43_sram;
wire [0:2] mux_tree_tapbuf_size6_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_44_sram;
wire [0:2] mux_tree_tapbuf_size6_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_45_sram;
wire [0:2] mux_tree_tapbuf_size6_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_46_sram;
wire [0:2] mux_tree_tapbuf_size6_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_47_sram;
wire [0:2] mux_tree_tapbuf_size6_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_48_sram;
wire [0:2] mux_tree_tapbuf_size6_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_49_sram;
wire [0:2] mux_tree_tapbuf_size6_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_50_sram;
wire [0:2] mux_tree_tapbuf_size6_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_51_sram;
wire [0:2] mux_tree_tapbuf_size6_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_52_sram;
wire [0:2] mux_tree_tapbuf_size6_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_53_sram;
wire [0:2] mux_tree_tapbuf_size6_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_54_sram;
wire [0:2] mux_tree_tapbuf_size6_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_55_sram;
wire [0:2] mux_tree_tapbuf_size6_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_56_sram;
wire [0:2] mux_tree_tapbuf_size6_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_57_sram;
wire [0:2] mux_tree_tapbuf_size6_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_58_sram;
wire [0:2] mux_tree_tapbuf_size6_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_59_sram;
wire [0:2] mux_tree_tapbuf_size6_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_60_sram;
wire [0:2] mux_tree_tapbuf_size6_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_61_sram;
wire [0:2] mux_tree_tapbuf_size6_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_62_sram;
wire [0:2] mux_tree_tapbuf_size6_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_63_sram;
wire [0:2] mux_tree_tapbuf_size6_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_64_sram;
wire [0:2] mux_tree_tapbuf_size6_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_65_sram;
wire [0:2] mux_tree_tapbuf_size6_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_66_sram;
wire [0:2] mux_tree_tapbuf_size6_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_67_sram;
wire [0:2] mux_tree_tapbuf_size6_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_68_sram;
wire [0:2] mux_tree_tapbuf_size6_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_69_sram;
wire [0:2] mux_tree_tapbuf_size6_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_70_sram;
wire [0:2] mux_tree_tapbuf_size6_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_71_sram;
wire [0:2] mux_tree_tapbuf_size6_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_72_sram;
wire [0:2] mux_tree_tapbuf_size6_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_73_sram;
wire [0:2] mux_tree_tapbuf_size6_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_74_sram;
wire [0:2] mux_tree_tapbuf_size6_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_75_sram;
wire [0:2] mux_tree_tapbuf_size6_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_76_sram;
wire [0:2] mux_tree_tapbuf_size6_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_77_sram;
wire [0:2] mux_tree_tapbuf_size6_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_78_sram;
wire [0:2] mux_tree_tapbuf_size6_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_79_sram;
wire [0:2] mux_tree_tapbuf_size6_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_80_sram;
wire [0:2] mux_tree_tapbuf_size6_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_81_sram;
wire [0:2] mux_tree_tapbuf_size6_81_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_82_sram;
wire [0:2] mux_tree_tapbuf_size6_82_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_83_sram;
wire [0:2] mux_tree_tapbuf_size6_83_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_84_sram;
wire [0:2] mux_tree_tapbuf_size6_84_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_85_sram;
wire [0:2] mux_tree_tapbuf_size6_85_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_86_sram;
wire [0:2] mux_tree_tapbuf_size6_86_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_87_sram;
wire [0:2] mux_tree_tapbuf_size6_87_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_88_sram;
wire [0:2] mux_tree_tapbuf_size6_88_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_89_sram;
wire [0:2] mux_tree_tapbuf_size6_89_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_90_sram;
wire [0:2] mux_tree_tapbuf_size6_90_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_91_sram;
wire [0:2] mux_tree_tapbuf_size6_91_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_92_sram;
wire [0:2] mux_tree_tapbuf_size6_92_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_93_sram;
wire [0:2] mux_tree_tapbuf_size6_93_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_94_sram;
wire [0:2] mux_tree_tapbuf_size6_94_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_95_sram;
wire [0:2] mux_tree_tapbuf_size6_95_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_96_sram;
wire [0:2] mux_tree_tapbuf_size6_96_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_97_sram;
wire [0:2] mux_tree_tapbuf_size6_97_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_98_sram;
wire [0:2] mux_tree_tapbuf_size6_98_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_99_sram;
wire [0:2] mux_tree_tapbuf_size6_99_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[177] = chanx_right_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[178] = chanx_right_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[179] = chanx_right_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[181] = chanx_right_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[182] = chanx_right_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[183] = chanx_right_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[185] = chanx_right_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[186] = chanx_right_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[187] = chanx_right_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[189] = chanx_right_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[190] = chanx_right_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[191] = chanx_right_in[190];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[193] = chanx_right_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[194] = chanx_right_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[195] = chanx_right_in[194];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[197] = chanx_right_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[198] = chanx_right_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[199] = chanx_right_in[198];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[201] = chanx_right_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[202] = chanx_right_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[203] = chanx_right_in[202];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[205] = chanx_right_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[206] = chanx_right_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[207] = chanx_right_in[206];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[209] = chanx_right_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[210] = chanx_right_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[211] = chanx_right_in[210];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[213] = chanx_right_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[214] = chanx_right_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[215] = chanx_right_in[214];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[217] = chanx_right_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[218] = chanx_right_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[219] = chanx_right_in[218];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[221] = chanx_right_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[222] = chanx_right_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[223] = chanx_right_in[222];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[225] = chanx_right_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[226] = chanx_right_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[227] = chanx_right_in[226];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[229] = chanx_right_in[228];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[230] = chanx_right_in[229];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[231] = chanx_right_in[230];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[233] = chanx_right_in[232];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[234] = chanx_right_in[233];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[235] = chanx_right_in[234];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[237] = chanx_right_in[236];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[238] = chanx_right_in[237];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[239] = chanx_right_in[238];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[241] = chanx_right_in[240];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[242] = chanx_right_in[241];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[243] = chanx_right_in[242];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[245] = chanx_right_in[244];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[246] = chanx_right_in[245];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[247] = chanx_right_in[246];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[249] = chanx_right_in[248];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[250] = chanx_right_in[249];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[251] = chanx_right_in[250];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[253] = chanx_right_in[252];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[254] = chanx_right_in[253];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[255] = chanx_right_in[254];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[257] = chanx_right_in[256];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[258] = chanx_right_in[257];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[259] = chanx_right_in[258];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[261] = chanx_right_in[260];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[262] = chanx_right_in[261];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[263] = chanx_right_in[262];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[265] = chanx_right_in[264];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[266] = chanx_right_in[265];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[267] = chanx_right_in[266];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[269] = chanx_right_in[268];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[270] = chanx_right_in[269];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[271] = chanx_right_in[270];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[273] = chanx_right_in[272];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[274] = chanx_right_in[273];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[275] = chanx_right_in[274];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[277] = chanx_right_in[276];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[278] = chanx_right_in[277];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[279] = chanx_right_in[278];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[281] = chanx_right_in[280];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[282] = chanx_right_in[281];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_left_out[283] = chanx_right_in[282];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 603 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 607 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 611 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 615 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 619 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 623 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 627 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 631 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 635 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 639 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 643 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 647 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 651 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 655 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 659 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 663 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 667 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 671 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 675 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 679 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 683 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 687 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 691 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 695 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 699 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 703 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 707 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 711 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 714 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 715 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 718 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 719 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 722 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 723 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 726 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 727 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 730 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 731 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 734 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 735 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 738 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 739 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 742 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 743 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 746 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 747 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 750 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 751 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 754 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 755 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 758 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 759 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 762 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 763 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 766 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 767 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 770 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 771 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 774 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 775 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- Local connection due to Wire 778 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[177] = chanx_left_in[176];
// ----- Local connection due to Wire 779 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[178] = chanx_left_in[177];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[179] = chanx_left_in[178];
// ----- Local connection due to Wire 782 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[181] = chanx_left_in[180];
// ----- Local connection due to Wire 783 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[182] = chanx_left_in[181];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[183] = chanx_left_in[182];
// ----- Local connection due to Wire 786 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[185] = chanx_left_in[184];
// ----- Local connection due to Wire 787 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[186] = chanx_left_in[185];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[187] = chanx_left_in[186];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[189] = chanx_left_in[188];
// ----- Local connection due to Wire 791 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[190] = chanx_left_in[189];
// ----- Local connection due to Wire 792 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[191] = chanx_left_in[190];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[193] = chanx_left_in[192];
// ----- Local connection due to Wire 795 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[194] = chanx_left_in[193];
// ----- Local connection due to Wire 796 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[195] = chanx_left_in[194];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[197] = chanx_left_in[196];
// ----- Local connection due to Wire 799 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[198] = chanx_left_in[197];
// ----- Local connection due to Wire 800 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[199] = chanx_left_in[198];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[201] = chanx_left_in[200];
// ----- Local connection due to Wire 803 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[202] = chanx_left_in[201];
// ----- Local connection due to Wire 804 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[203] = chanx_left_in[202];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[205] = chanx_left_in[204];
// ----- Local connection due to Wire 807 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[206] = chanx_left_in[205];
// ----- Local connection due to Wire 808 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[207] = chanx_left_in[206];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[209] = chanx_left_in[208];
// ----- Local connection due to Wire 811 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[210] = chanx_left_in[209];
// ----- Local connection due to Wire 812 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[211] = chanx_left_in[210];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[213] = chanx_left_in[212];
// ----- Local connection due to Wire 815 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[214] = chanx_left_in[213];
// ----- Local connection due to Wire 816 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[215] = chanx_left_in[214];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[217] = chanx_left_in[216];
// ----- Local connection due to Wire 819 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[218] = chanx_left_in[217];
// ----- Local connection due to Wire 820 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[219] = chanx_left_in[218];
// ----- Local connection due to Wire 822 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[221] = chanx_left_in[220];
// ----- Local connection due to Wire 823 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[222] = chanx_left_in[221];
// ----- Local connection due to Wire 824 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[223] = chanx_left_in[222];
// ----- Local connection due to Wire 826 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[225] = chanx_left_in[224];
// ----- Local connection due to Wire 827 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[226] = chanx_left_in[225];
// ----- Local connection due to Wire 828 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[227] = chanx_left_in[226];
// ----- Local connection due to Wire 830 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[229] = chanx_left_in[228];
// ----- Local connection due to Wire 831 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[230] = chanx_left_in[229];
// ----- Local connection due to Wire 832 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[231] = chanx_left_in[230];
// ----- Local connection due to Wire 834 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[233] = chanx_left_in[232];
// ----- Local connection due to Wire 835 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[234] = chanx_left_in[233];
// ----- Local connection due to Wire 836 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[235] = chanx_left_in[234];
// ----- Local connection due to Wire 838 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[237] = chanx_left_in[236];
// ----- Local connection due to Wire 839 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[238] = chanx_left_in[237];
// ----- Local connection due to Wire 840 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[239] = chanx_left_in[238];
// ----- Local connection due to Wire 842 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[241] = chanx_left_in[240];
// ----- Local connection due to Wire 843 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[242] = chanx_left_in[241];
// ----- Local connection due to Wire 844 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[243] = chanx_left_in[242];
// ----- Local connection due to Wire 846 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[245] = chanx_left_in[244];
// ----- Local connection due to Wire 847 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[246] = chanx_left_in[245];
// ----- Local connection due to Wire 848 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[247] = chanx_left_in[246];
// ----- Local connection due to Wire 850 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[249] = chanx_left_in[248];
// ----- Local connection due to Wire 851 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[250] = chanx_left_in[249];
// ----- Local connection due to Wire 852 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[251] = chanx_left_in[250];
// ----- Local connection due to Wire 854 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[253] = chanx_left_in[252];
// ----- Local connection due to Wire 855 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[254] = chanx_left_in[253];
// ----- Local connection due to Wire 856 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[255] = chanx_left_in[254];
// ----- Local connection due to Wire 858 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[257] = chanx_left_in[256];
// ----- Local connection due to Wire 859 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[258] = chanx_left_in[257];
// ----- Local connection due to Wire 860 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[259] = chanx_left_in[258];
// ----- Local connection due to Wire 862 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[261] = chanx_left_in[260];
// ----- Local connection due to Wire 863 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[262] = chanx_left_in[261];
// ----- Local connection due to Wire 864 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[263] = chanx_left_in[262];
// ----- Local connection due to Wire 866 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[265] = chanx_left_in[264];
// ----- Local connection due to Wire 867 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[266] = chanx_left_in[265];
// ----- Local connection due to Wire 868 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[267] = chanx_left_in[266];
// ----- Local connection due to Wire 870 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[269] = chanx_left_in[268];
// ----- Local connection due to Wire 871 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[270] = chanx_left_in[269];
// ----- Local connection due to Wire 872 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[271] = chanx_left_in[270];
// ----- Local connection due to Wire 874 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[273] = chanx_left_in[272];
// ----- Local connection due to Wire 875 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[274] = chanx_left_in[273];
// ----- Local connection due to Wire 876 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[275] = chanx_left_in[274];
// ----- Local connection due to Wire 878 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[277] = chanx_left_in[276];
// ----- Local connection due to Wire 879 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[278] = chanx_left_in[277];
// ----- Local connection due to Wire 880 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[279] = chanx_left_in[278];
// ----- Local connection due to Wire 882 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[281] = chanx_left_in[280];
// ----- Local connection due to Wire 883 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[282] = chanx_left_in[281];
// ----- Local connection due to Wire 884 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chanx_right_out[283] = chanx_left_in[282];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size5 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[70], chany_bottom_in[142], chany_bottom_in[214]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size5 mux_right_track_8 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[69], chany_bottom_in[141], chany_bottom_in[213]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size5 mux_right_track_56 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[63], chany_bottom_in[135], chany_bottom_in[207], chany_bottom_in[279]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size5 mux_right_track_64 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[62], chany_bottom_in[134], chany_bottom_in[206], chany_bottom_in[278]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size5 mux_right_track_128 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[54], chany_bottom_in[126], chany_bottom_in[198], chany_bottom_in[270]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size5 mux_right_track_136 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[53], chany_bottom_in[125], chany_bottom_in[197], chany_bottom_in[269]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size5 mux_right_track_200 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[45], chany_bottom_in[117], chany_bottom_in[189], chany_bottom_in[261]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size5 mux_right_track_208 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[44], chany_bottom_in[116], chany_bottom_in[188], chany_bottom_in[260]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size5 mux_right_track_272 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[36], chany_bottom_in[108], chany_bottom_in[180], chany_bottom_in[252]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size5 mux_right_track_280 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[35], chany_bottom_in[107], chany_bottom_in[179], chany_bottom_in[251]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size5 mux_right_track_344 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[27], chany_bottom_in[99], chany_bottom_in[171], chany_bottom_in[243]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size5 mux_right_track_352 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[26], chany_bottom_in[98], chany_bottom_in[170], chany_bottom_in[242]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size5 mux_right_track_416 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[18], chany_bottom_in[90], chany_bottom_in[162], chany_bottom_in[234]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chanx_right_out[208]));

	mux_tree_tapbuf_size5 mux_right_track_424 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[17], chany_bottom_in[89], chany_bottom_in[161], chany_bottom_in[233]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chanx_right_out[212]));

	mux_tree_tapbuf_size5 mux_right_track_488 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[9], chany_bottom_in[81], chany_bottom_in[153], chany_bottom_in[225]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chanx_right_out[244]));

	mux_tree_tapbuf_size5 mux_right_track_496 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[8], chany_bottom_in[80], chany_bottom_in[152], chany_bottom_in[224]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chanx_right_out[248]));

	mux_tree_tapbuf_size5 mux_right_track_560 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[0], chany_bottom_in[72], chany_bottom_in[144], chany_bottom_in[216]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chanx_right_out[280]));

	mux_tree_tapbuf_size5 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[1], chanx_left_in[7]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size5 mux_bottom_track_19 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[13], chanx_left_in[43]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_bottom_out[9]));

	mux_tree_tapbuf_size5 mux_left_track_1 (
		.in({chany_bottom_in[71], chany_bottom_in[143], chany_bottom_in[215], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size5 mux_left_track_57 (
		.in({chany_bottom_in[6], chany_bottom_in[78], chany_bottom_in[150], chany_bottom_in[222], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size5 mux_left_track_65 (
		.in({chany_bottom_in[7], chany_bottom_in[79], chany_bottom_in[151], chany_bottom_in[223], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size5 mux_left_track_129 (
		.in({chany_bottom_in[15], chany_bottom_in[87], chany_bottom_in[159], chany_bottom_in[231], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size5 mux_left_track_137 (
		.in({chany_bottom_in[16], chany_bottom_in[88], chany_bottom_in[160], chany_bottom_in[232], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size5 mux_left_track_201 (
		.in({chany_bottom_in[24], chany_bottom_in[96], chany_bottom_in[168], chany_bottom_in[240], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size5 mux_left_track_209 (
		.in({chany_bottom_in[25], chany_bottom_in[97], chany_bottom_in[169], chany_bottom_in[241], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size5 mux_left_track_273 (
		.in({chany_bottom_in[33], chany_bottom_in[105], chany_bottom_in[177], chany_bottom_in[249], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size5 mux_left_track_281 (
		.in({chany_bottom_in[34], chany_bottom_in[106], chany_bottom_in[178], chany_bottom_in[250], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size5 mux_left_track_345 (
		.in({chany_bottom_in[42], chany_bottom_in[114], chany_bottom_in[186], chany_bottom_in[258], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size5 mux_left_track_353 (
		.in({chany_bottom_in[43], chany_bottom_in[115], chany_bottom_in[187], chany_bottom_in[259], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size5 mux_left_track_417 (
		.in({chany_bottom_in[51], chany_bottom_in[123], chany_bottom_in[195], chany_bottom_in[267], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chanx_left_out[208]));

	mux_tree_tapbuf_size5 mux_left_track_425 (
		.in({chany_bottom_in[52], chany_bottom_in[124], chany_bottom_in[196], chany_bottom_in[268], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chanx_left_out[212]));

	mux_tree_tapbuf_size5 mux_left_track_489 (
		.in({chany_bottom_in[60], chany_bottom_in[132], chany_bottom_in[204], chany_bottom_in[276], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chanx_left_out[244]));

	mux_tree_tapbuf_size5 mux_left_track_497 (
		.in({chany_bottom_in[61], chany_bottom_in[133], chany_bottom_in[205], chany_bottom_in[277], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chanx_left_out[248]));

	mux_tree_tapbuf_size5_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_right_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_left_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_right_track_16 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[68], chany_bottom_in[140], chany_bottom_in[212], chany_bottom_in[284]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size6 mux_right_track_24 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[67], chany_bottom_in[139], chany_bottom_in[211], chany_bottom_in[283]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size6 mux_right_track_32 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[66], chany_bottom_in[138], chany_bottom_in[210], chany_bottom_in[282]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size6 mux_right_track_40 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[65], chany_bottom_in[137], chany_bottom_in[209], chany_bottom_in[281]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size6 mux_right_track_48 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[64], chany_bottom_in[136], chany_bottom_in[208], chany_bottom_in[280]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size6 mux_right_track_72 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[61], chany_bottom_in[133], chany_bottom_in[205], chany_bottom_in[277]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size6 mux_right_track_80 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[60], chany_bottom_in[132], chany_bottom_in[204], chany_bottom_in[276]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size6 mux_right_track_88 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[59], chany_bottom_in[131], chany_bottom_in[203], chany_bottom_in[275]}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size6 mux_right_track_96 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[58], chany_bottom_in[130], chany_bottom_in[202], chany_bottom_in[274]}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size6 mux_right_track_104 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[57], chany_bottom_in[129], chany_bottom_in[201], chany_bottom_in[273]}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size6 mux_right_track_112 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[56], chany_bottom_in[128], chany_bottom_in[200], chany_bottom_in[272]}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size6 mux_right_track_120 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[55], chany_bottom_in[127], chany_bottom_in[199], chany_bottom_in[271]}),
		.sram(mux_tree_tapbuf_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_11_sram_inv[0:2]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size6 mux_right_track_144 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[52], chany_bottom_in[124], chany_bottom_in[196], chany_bottom_in[268]}),
		.sram(mux_tree_tapbuf_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_12_sram_inv[0:2]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size6 mux_right_track_152 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[51], chany_bottom_in[123], chany_bottom_in[195], chany_bottom_in[267]}),
		.sram(mux_tree_tapbuf_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_13_sram_inv[0:2]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size6 mux_right_track_160 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[50], chany_bottom_in[122], chany_bottom_in[194], chany_bottom_in[266]}),
		.sram(mux_tree_tapbuf_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_14_sram_inv[0:2]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size6 mux_right_track_168 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[49], chany_bottom_in[121], chany_bottom_in[193], chany_bottom_in[265]}),
		.sram(mux_tree_tapbuf_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_15_sram_inv[0:2]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size6 mux_right_track_176 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[48], chany_bottom_in[120], chany_bottom_in[192], chany_bottom_in[264]}),
		.sram(mux_tree_tapbuf_size6_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_16_sram_inv[0:2]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size6 mux_right_track_184 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[47], chany_bottom_in[119], chany_bottom_in[191], chany_bottom_in[263]}),
		.sram(mux_tree_tapbuf_size6_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_17_sram_inv[0:2]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size6 mux_right_track_192 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[46], chany_bottom_in[118], chany_bottom_in[190], chany_bottom_in[262]}),
		.sram(mux_tree_tapbuf_size6_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_18_sram_inv[0:2]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size6 mux_right_track_216 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[43], chany_bottom_in[115], chany_bottom_in[187], chany_bottom_in[259]}),
		.sram(mux_tree_tapbuf_size6_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_19_sram_inv[0:2]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size6 mux_right_track_224 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[42], chany_bottom_in[114], chany_bottom_in[186], chany_bottom_in[258]}),
		.sram(mux_tree_tapbuf_size6_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_20_sram_inv[0:2]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size6 mux_right_track_232 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[41], chany_bottom_in[113], chany_bottom_in[185], chany_bottom_in[257]}),
		.sram(mux_tree_tapbuf_size6_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_21_sram_inv[0:2]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size6 mux_right_track_240 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[40], chany_bottom_in[112], chany_bottom_in[184], chany_bottom_in[256]}),
		.sram(mux_tree_tapbuf_size6_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_22_sram_inv[0:2]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size6 mux_right_track_248 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[39], chany_bottom_in[111], chany_bottom_in[183], chany_bottom_in[255]}),
		.sram(mux_tree_tapbuf_size6_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_23_sram_inv[0:2]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size6 mux_right_track_256 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[38], chany_bottom_in[110], chany_bottom_in[182], chany_bottom_in[254]}),
		.sram(mux_tree_tapbuf_size6_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_24_sram_inv[0:2]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size6 mux_right_track_264 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[37], chany_bottom_in[109], chany_bottom_in[181], chany_bottom_in[253]}),
		.sram(mux_tree_tapbuf_size6_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_25_sram_inv[0:2]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size6 mux_right_track_288 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[34], chany_bottom_in[106], chany_bottom_in[178], chany_bottom_in[250]}),
		.sram(mux_tree_tapbuf_size6_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_26_sram_inv[0:2]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size6 mux_right_track_296 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[33], chany_bottom_in[105], chany_bottom_in[177], chany_bottom_in[249]}),
		.sram(mux_tree_tapbuf_size6_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_27_sram_inv[0:2]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size6 mux_right_track_304 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[32], chany_bottom_in[104], chany_bottom_in[176], chany_bottom_in[248]}),
		.sram(mux_tree_tapbuf_size6_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_28_sram_inv[0:2]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size6 mux_right_track_312 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[31], chany_bottom_in[103], chany_bottom_in[175], chany_bottom_in[247]}),
		.sram(mux_tree_tapbuf_size6_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_29_sram_inv[0:2]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size6 mux_right_track_320 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[30], chany_bottom_in[102], chany_bottom_in[174], chany_bottom_in[246]}),
		.sram(mux_tree_tapbuf_size6_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_30_sram_inv[0:2]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size6 mux_right_track_328 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[29], chany_bottom_in[101], chany_bottom_in[173], chany_bottom_in[245]}),
		.sram(mux_tree_tapbuf_size6_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_31_sram_inv[0:2]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size6 mux_right_track_336 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[28], chany_bottom_in[100], chany_bottom_in[172], chany_bottom_in[244]}),
		.sram(mux_tree_tapbuf_size6_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_32_sram_inv[0:2]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size6 mux_right_track_360 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[25], chany_bottom_in[97], chany_bottom_in[169], chany_bottom_in[241]}),
		.sram(mux_tree_tapbuf_size6_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_33_sram_inv[0:2]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size6 mux_right_track_368 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[24], chany_bottom_in[96], chany_bottom_in[168], chany_bottom_in[240]}),
		.sram(mux_tree_tapbuf_size6_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_34_sram_inv[0:2]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size6 mux_right_track_376 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[23], chany_bottom_in[95], chany_bottom_in[167], chany_bottom_in[239]}),
		.sram(mux_tree_tapbuf_size6_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_35_sram_inv[0:2]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size6 mux_right_track_384 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[22], chany_bottom_in[94], chany_bottom_in[166], chany_bottom_in[238]}),
		.sram(mux_tree_tapbuf_size6_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_36_sram_inv[0:2]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size6 mux_right_track_392 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[21], chany_bottom_in[93], chany_bottom_in[165], chany_bottom_in[237]}),
		.sram(mux_tree_tapbuf_size6_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_37_sram_inv[0:2]),
		.out(chanx_right_out[196]));

	mux_tree_tapbuf_size6 mux_right_track_400 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[20], chany_bottom_in[92], chany_bottom_in[164], chany_bottom_in[236]}),
		.sram(mux_tree_tapbuf_size6_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_38_sram_inv[0:2]),
		.out(chanx_right_out[200]));

	mux_tree_tapbuf_size6 mux_right_track_408 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[19], chany_bottom_in[91], chany_bottom_in[163], chany_bottom_in[235]}),
		.sram(mux_tree_tapbuf_size6_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_39_sram_inv[0:2]),
		.out(chanx_right_out[204]));

	mux_tree_tapbuf_size6 mux_right_track_432 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[16], chany_bottom_in[88], chany_bottom_in[160], chany_bottom_in[232]}),
		.sram(mux_tree_tapbuf_size6_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_40_sram_inv[0:2]),
		.out(chanx_right_out[216]));

	mux_tree_tapbuf_size6 mux_right_track_440 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[15], chany_bottom_in[87], chany_bottom_in[159], chany_bottom_in[231]}),
		.sram(mux_tree_tapbuf_size6_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_41_sram_inv[0:2]),
		.out(chanx_right_out[220]));

	mux_tree_tapbuf_size6 mux_right_track_448 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[14], chany_bottom_in[86], chany_bottom_in[158], chany_bottom_in[230]}),
		.sram(mux_tree_tapbuf_size6_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_42_sram_inv[0:2]),
		.out(chanx_right_out[224]));

	mux_tree_tapbuf_size6 mux_right_track_456 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[13], chany_bottom_in[85], chany_bottom_in[157], chany_bottom_in[229]}),
		.sram(mux_tree_tapbuf_size6_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_43_sram_inv[0:2]),
		.out(chanx_right_out[228]));

	mux_tree_tapbuf_size6 mux_right_track_464 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[12], chany_bottom_in[84], chany_bottom_in[156], chany_bottom_in[228]}),
		.sram(mux_tree_tapbuf_size6_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_44_sram_inv[0:2]),
		.out(chanx_right_out[232]));

	mux_tree_tapbuf_size6 mux_right_track_472 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[11], chany_bottom_in[83], chany_bottom_in[155], chany_bottom_in[227]}),
		.sram(mux_tree_tapbuf_size6_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_45_sram_inv[0:2]),
		.out(chanx_right_out[236]));

	mux_tree_tapbuf_size6 mux_right_track_480 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[10], chany_bottom_in[82], chany_bottom_in[154], chany_bottom_in[226]}),
		.sram(mux_tree_tapbuf_size6_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_46_sram_inv[0:2]),
		.out(chanx_right_out[240]));

	mux_tree_tapbuf_size6 mux_right_track_504 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[7], chany_bottom_in[79], chany_bottom_in[151], chany_bottom_in[223]}),
		.sram(mux_tree_tapbuf_size6_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_47_sram_inv[0:2]),
		.out(chanx_right_out[252]));

	mux_tree_tapbuf_size6 mux_right_track_512 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[6], chany_bottom_in[78], chany_bottom_in[150], chany_bottom_in[222]}),
		.sram(mux_tree_tapbuf_size6_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_48_sram_inv[0:2]),
		.out(chanx_right_out[256]));

	mux_tree_tapbuf_size6 mux_right_track_520 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[5], chany_bottom_in[77], chany_bottom_in[149], chany_bottom_in[221]}),
		.sram(mux_tree_tapbuf_size6_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_49_sram_inv[0:2]),
		.out(chanx_right_out[260]));

	mux_tree_tapbuf_size6 mux_right_track_528 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[4], chany_bottom_in[76], chany_bottom_in[148], chany_bottom_in[220]}),
		.sram(mux_tree_tapbuf_size6_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_50_sram_inv[0:2]),
		.out(chanx_right_out[264]));

	mux_tree_tapbuf_size6 mux_right_track_536 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[3], chany_bottom_in[75], chany_bottom_in[147], chany_bottom_in[219]}),
		.sram(mux_tree_tapbuf_size6_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_51_sram_inv[0:2]),
		.out(chanx_right_out[268]));

	mux_tree_tapbuf_size6 mux_right_track_544 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[2], chany_bottom_in[74], chany_bottom_in[146], chany_bottom_in[218]}),
		.sram(mux_tree_tapbuf_size6_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_52_sram_inv[0:2]),
		.out(chanx_right_out[272]));

	mux_tree_tapbuf_size6 mux_right_track_552 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[1], chany_bottom_in[73], chany_bottom_in[145], chany_bottom_in[217]}),
		.sram(mux_tree_tapbuf_size6_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_53_sram_inv[0:2]),
		.out(chanx_right_out[276]));

	mux_tree_tapbuf_size6 mux_left_track_9 (
		.in({chany_bottom_in[0], chany_bottom_in[72], chany_bottom_in[144], chany_bottom_in[216], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_54_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size6 mux_left_track_17 (
		.in({chany_bottom_in[1], chany_bottom_in[73], chany_bottom_in[145], chany_bottom_in[217], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_55_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size6 mux_left_track_25 (
		.in({chany_bottom_in[2], chany_bottom_in[74], chany_bottom_in[146], chany_bottom_in[218], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_56_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size6 mux_left_track_33 (
		.in({chany_bottom_in[3], chany_bottom_in[75], chany_bottom_in[147], chany_bottom_in[219], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_57_sram_inv[0:2]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size6 mux_left_track_41 (
		.in({chany_bottom_in[4], chany_bottom_in[76], chany_bottom_in[148], chany_bottom_in[220], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_58_sram_inv[0:2]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size6 mux_left_track_49 (
		.in({chany_bottom_in[5], chany_bottom_in[77], chany_bottom_in[149], chany_bottom_in[221], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_59_sram_inv[0:2]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size6 mux_left_track_73 (
		.in({chany_bottom_in[8], chany_bottom_in[80], chany_bottom_in[152], chany_bottom_in[224], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_60_sram_inv[0:2]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size6 mux_left_track_81 (
		.in({chany_bottom_in[9], chany_bottom_in[81], chany_bottom_in[153], chany_bottom_in[225], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_61_sram_inv[0:2]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size6 mux_left_track_89 (
		.in({chany_bottom_in[10], chany_bottom_in[82], chany_bottom_in[154], chany_bottom_in[226], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_62_sram_inv[0:2]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size6 mux_left_track_97 (
		.in({chany_bottom_in[11], chany_bottom_in[83], chany_bottom_in[155], chany_bottom_in[227], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_63_sram_inv[0:2]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size6 mux_left_track_105 (
		.in({chany_bottom_in[12], chany_bottom_in[84], chany_bottom_in[156], chany_bottom_in[228], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_64_sram_inv[0:2]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size6 mux_left_track_113 (
		.in({chany_bottom_in[13], chany_bottom_in[85], chany_bottom_in[157], chany_bottom_in[229], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_65_sram_inv[0:2]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size6 mux_left_track_121 (
		.in({chany_bottom_in[14], chany_bottom_in[86], chany_bottom_in[158], chany_bottom_in[230], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_66_sram_inv[0:2]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size6 mux_left_track_145 (
		.in({chany_bottom_in[17], chany_bottom_in[89], chany_bottom_in[161], chany_bottom_in[233], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_67_sram_inv[0:2]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size6 mux_left_track_153 (
		.in({chany_bottom_in[18], chany_bottom_in[90], chany_bottom_in[162], chany_bottom_in[234], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_68_sram_inv[0:2]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size6 mux_left_track_161 (
		.in({chany_bottom_in[19], chany_bottom_in[91], chany_bottom_in[163], chany_bottom_in[235], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_69_sram_inv[0:2]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size6 mux_left_track_169 (
		.in({chany_bottom_in[20], chany_bottom_in[92], chany_bottom_in[164], chany_bottom_in[236], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_70_sram_inv[0:2]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size6 mux_left_track_177 (
		.in({chany_bottom_in[21], chany_bottom_in[93], chany_bottom_in[165], chany_bottom_in[237], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_71_sram_inv[0:2]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size6 mux_left_track_185 (
		.in({chany_bottom_in[22], chany_bottom_in[94], chany_bottom_in[166], chany_bottom_in[238], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_72_sram_inv[0:2]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size6 mux_left_track_193 (
		.in({chany_bottom_in[23], chany_bottom_in[95], chany_bottom_in[167], chany_bottom_in[239], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_73_sram_inv[0:2]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size6 mux_left_track_217 (
		.in({chany_bottom_in[26], chany_bottom_in[98], chany_bottom_in[170], chany_bottom_in[242], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_74_sram_inv[0:2]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size6 mux_left_track_225 (
		.in({chany_bottom_in[27], chany_bottom_in[99], chany_bottom_in[171], chany_bottom_in[243], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_75_sram_inv[0:2]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size6 mux_left_track_233 (
		.in({chany_bottom_in[28], chany_bottom_in[100], chany_bottom_in[172], chany_bottom_in[244], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_76_sram_inv[0:2]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size6 mux_left_track_241 (
		.in({chany_bottom_in[29], chany_bottom_in[101], chany_bottom_in[173], chany_bottom_in[245], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_77_sram_inv[0:2]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size6 mux_left_track_249 (
		.in({chany_bottom_in[30], chany_bottom_in[102], chany_bottom_in[174], chany_bottom_in[246], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_78_sram_inv[0:2]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size6 mux_left_track_257 (
		.in({chany_bottom_in[31], chany_bottom_in[103], chany_bottom_in[175], chany_bottom_in[247], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_79_sram_inv[0:2]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size6 mux_left_track_265 (
		.in({chany_bottom_in[32], chany_bottom_in[104], chany_bottom_in[176], chany_bottom_in[248], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_80_sram_inv[0:2]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size6 mux_left_track_289 (
		.in({chany_bottom_in[35], chany_bottom_in[107], chany_bottom_in[179], chany_bottom_in[251], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_81_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_81_sram_inv[0:2]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size6 mux_left_track_297 (
		.in({chany_bottom_in[36], chany_bottom_in[108], chany_bottom_in[180], chany_bottom_in[252], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_82_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_82_sram_inv[0:2]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size6 mux_left_track_305 (
		.in({chany_bottom_in[37], chany_bottom_in[109], chany_bottom_in[181], chany_bottom_in[253], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_83_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_83_sram_inv[0:2]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size6 mux_left_track_313 (
		.in({chany_bottom_in[38], chany_bottom_in[110], chany_bottom_in[182], chany_bottom_in[254], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_84_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_84_sram_inv[0:2]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size6 mux_left_track_321 (
		.in({chany_bottom_in[39], chany_bottom_in[111], chany_bottom_in[183], chany_bottom_in[255], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_85_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_85_sram_inv[0:2]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size6 mux_left_track_329 (
		.in({chany_bottom_in[40], chany_bottom_in[112], chany_bottom_in[184], chany_bottom_in[256], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_86_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_86_sram_inv[0:2]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size6 mux_left_track_337 (
		.in({chany_bottom_in[41], chany_bottom_in[113], chany_bottom_in[185], chany_bottom_in[257], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_87_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_87_sram_inv[0:2]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size6 mux_left_track_361 (
		.in({chany_bottom_in[44], chany_bottom_in[116], chany_bottom_in[188], chany_bottom_in[260], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_88_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_88_sram_inv[0:2]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size6 mux_left_track_369 (
		.in({chany_bottom_in[45], chany_bottom_in[117], chany_bottom_in[189], chany_bottom_in[261], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_89_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_89_sram_inv[0:2]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size6 mux_left_track_377 (
		.in({chany_bottom_in[46], chany_bottom_in[118], chany_bottom_in[190], chany_bottom_in[262], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_90_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_90_sram_inv[0:2]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size6 mux_left_track_385 (
		.in({chany_bottom_in[47], chany_bottom_in[119], chany_bottom_in[191], chany_bottom_in[263], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_91_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_91_sram_inv[0:2]),
		.out(chanx_left_out[192]));

	mux_tree_tapbuf_size6 mux_left_track_393 (
		.in({chany_bottom_in[48], chany_bottom_in[120], chany_bottom_in[192], chany_bottom_in[264], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_92_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_92_sram_inv[0:2]),
		.out(chanx_left_out[196]));

	mux_tree_tapbuf_size6 mux_left_track_401 (
		.in({chany_bottom_in[49], chany_bottom_in[121], chany_bottom_in[193], chany_bottom_in[265], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_93_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_93_sram_inv[0:2]),
		.out(chanx_left_out[200]));

	mux_tree_tapbuf_size6 mux_left_track_409 (
		.in({chany_bottom_in[50], chany_bottom_in[122], chany_bottom_in[194], chany_bottom_in[266], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_94_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_94_sram_inv[0:2]),
		.out(chanx_left_out[204]));

	mux_tree_tapbuf_size6 mux_left_track_433 (
		.in({chany_bottom_in[53], chany_bottom_in[125], chany_bottom_in[197], chany_bottom_in[269], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_95_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_95_sram_inv[0:2]),
		.out(chanx_left_out[216]));

	mux_tree_tapbuf_size6 mux_left_track_441 (
		.in({chany_bottom_in[54], chany_bottom_in[126], chany_bottom_in[198], chany_bottom_in[270], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_96_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_96_sram_inv[0:2]),
		.out(chanx_left_out[220]));

	mux_tree_tapbuf_size6 mux_left_track_449 (
		.in({chany_bottom_in[55], chany_bottom_in[127], chany_bottom_in[199], chany_bottom_in[271], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_97_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_97_sram_inv[0:2]),
		.out(chanx_left_out[224]));

	mux_tree_tapbuf_size6 mux_left_track_457 (
		.in({chany_bottom_in[56], chany_bottom_in[128], chany_bottom_in[200], chany_bottom_in[272], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_98_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_98_sram_inv[0:2]),
		.out(chanx_left_out[228]));

	mux_tree_tapbuf_size6 mux_left_track_465 (
		.in({chany_bottom_in[57], chany_bottom_in[129], chany_bottom_in[201], chany_bottom_in[273], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_99_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_99_sram_inv[0:2]),
		.out(chanx_left_out[232]));

	mux_tree_tapbuf_size6 mux_left_track_473 (
		.in({chany_bottom_in[58], chany_bottom_in[130], chany_bottom_in[202], chany_bottom_in[274], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_100_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_100_sram_inv[0:2]),
		.out(chanx_left_out[236]));

	mux_tree_tapbuf_size6 mux_left_track_481 (
		.in({chany_bottom_in[59], chany_bottom_in[131], chany_bottom_in[203], chany_bottom_in[275], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_101_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_101_sram_inv[0:2]),
		.out(chanx_left_out[240]));

	mux_tree_tapbuf_size6 mux_left_track_505 (
		.in({chany_bottom_in[62], chany_bottom_in[134], chany_bottom_in[206], chany_bottom_in[278], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_102_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_102_sram_inv[0:2]),
		.out(chanx_left_out[252]));

	mux_tree_tapbuf_size6 mux_left_track_513 (
		.in({chany_bottom_in[63], chany_bottom_in[135], chany_bottom_in[207], chany_bottom_in[279], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_103_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_103_sram_inv[0:2]),
		.out(chanx_left_out[256]));

	mux_tree_tapbuf_size6 mux_left_track_521 (
		.in({chany_bottom_in[64], chany_bottom_in[136], chany_bottom_in[208], chany_bottom_in[280], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_104_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_104_sram_inv[0:2]),
		.out(chanx_left_out[260]));

	mux_tree_tapbuf_size6 mux_left_track_529 (
		.in({chany_bottom_in[65], chany_bottom_in[137], chany_bottom_in[209], chany_bottom_in[281], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_105_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_105_sram_inv[0:2]),
		.out(chanx_left_out[264]));

	mux_tree_tapbuf_size6 mux_left_track_537 (
		.in({chany_bottom_in[66], chany_bottom_in[138], chany_bottom_in[210], chany_bottom_in[282], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_106_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_106_sram_inv[0:2]),
		.out(chanx_left_out[268]));

	mux_tree_tapbuf_size6 mux_left_track_545 (
		.in({chany_bottom_in[67], chany_bottom_in[139], chany_bottom_in[211], chany_bottom_in[283], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_107_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_107_sram_inv[0:2]),
		.out(chanx_left_out[272]));

	mux_tree_tapbuf_size6 mux_left_track_553 (
		.in({chany_bottom_in[68], chany_bottom_in[140], chany_bottom_in[212], chany_bottom_in[284], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_108_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_108_sram_inv[0:2]),
		.out(chanx_left_out[276]));

	mux_tree_tapbuf_size6_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_16_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_17_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_18_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_19_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_20_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_21_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_22_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_23_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_24_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_25_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_26_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_27_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_28_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_29_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_30_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_31_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_32_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_33_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_34_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_35_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_36_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_37_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_38_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_39_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_40_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_41_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_42_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_43_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_44_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_45_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_46_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_47_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_48_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_49_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_50_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_51_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_52_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_right_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_53_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_54_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_55_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_56_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_57_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_58_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_59_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_60_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_61_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_62_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_63_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_64_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_65_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_66_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_67_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_68_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_69_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_70_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_71_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_72_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_73_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_74_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_75_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_76_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_77_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_78_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_79_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_80_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_81_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_81_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_82_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_82_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_83_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_83_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_84_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_84_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_85_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_85_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_86_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_86_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_87_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_87_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_88_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_88_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_89_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_89_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_90_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_90_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_91_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_91_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_92_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_92_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_93_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_93_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_94_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_94_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_95_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_95_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_96_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_96_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_97_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_97_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_98_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_98_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_99_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_99_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_100_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_100_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_101_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_101_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_102_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_102_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_103_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_103_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_104_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_104_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_105_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_105_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_106_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_106_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_107_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_107_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_left_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_108_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_108_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_right_track_568 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[71], chany_bottom_in[143], chany_bottom_in[215]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chanx_right_out[284]));

	mux_tree_tapbuf_size4 mux_bottom_track_3 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[2], chanx_left_in[11]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_bottom_out[1]));

	mux_tree_tapbuf_size4 mux_bottom_track_5 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[4], chanx_left_in[15]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_bottom_out[2]));

	mux_tree_tapbuf_size4 mux_bottom_track_7 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[5], chanx_left_in[19]}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chany_bottom_out[3]));

	mux_tree_tapbuf_size4 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[6], chanx_left_in[23]}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size4 mux_bottom_track_11 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[8], chanx_left_in[27]}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chany_bottom_out[5]));

	mux_tree_tapbuf_size4 mux_bottom_track_13 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[9], chanx_left_in[31]}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chany_bottom_out[6]));

	mux_tree_tapbuf_size4 mux_bottom_track_15 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[10], chanx_left_in[35]}),
		.sram(mux_tree_tapbuf_size4_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_7_sram_inv[0:2]),
		.out(chany_bottom_out[7]));

	mux_tree_tapbuf_size4 mux_bottom_track_17 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[12], chanx_left_in[39]}),
		.sram(mux_tree_tapbuf_size4_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_8_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size4 mux_bottom_track_21 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[14], chanx_left_in[47]}),
		.sram(mux_tree_tapbuf_size4_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_9_sram_inv[0:2]),
		.out(chany_bottom_out[10]));

	mux_tree_tapbuf_size4 mux_bottom_track_23 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[16], chanx_left_in[51]}),
		.sram(mux_tree_tapbuf_size4_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_10_sram_inv[0:2]),
		.out(chany_bottom_out[11]));

	mux_tree_tapbuf_size4 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[17], chanx_left_in[55]}),
		.sram(mux_tree_tapbuf_size4_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_11_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size4 mux_bottom_track_27 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[18], chanx_left_in[59]}),
		.sram(mux_tree_tapbuf_size4_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_12_sram_inv[0:2]),
		.out(chany_bottom_out[13]));

	mux_tree_tapbuf_size4 mux_bottom_track_29 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[20], chanx_left_in[63]}),
		.sram(mux_tree_tapbuf_size4_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_13_sram_inv[0:2]),
		.out(chany_bottom_out[14]));

	mux_tree_tapbuf_size4 mux_bottom_track_31 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[21], chanx_left_in[67]}),
		.sram(mux_tree_tapbuf_size4_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_14_sram_inv[0:2]),
		.out(chany_bottom_out[15]));

	mux_tree_tapbuf_size4 mux_bottom_track_37 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[25], chanx_left_in[79]}),
		.sram(mux_tree_tapbuf_size4_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_15_sram_inv[0:2]),
		.out(chany_bottom_out[18]));

	mux_tree_tapbuf_size4 mux_bottom_track_39 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[26], chanx_left_in[83]}),
		.sram(mux_tree_tapbuf_size4_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_16_sram_inv[0:2]),
		.out(chany_bottom_out[19]));

	mux_tree_tapbuf_size4 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[28], chanx_left_in[87]}),
		.sram(mux_tree_tapbuf_size4_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_17_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size4 mux_bottom_track_43 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[29], chanx_left_in[91]}),
		.sram(mux_tree_tapbuf_size4_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_18_sram_inv[0:2]),
		.out(chany_bottom_out[21]));

	mux_tree_tapbuf_size4 mux_bottom_track_45 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[30], chanx_left_in[95]}),
		.sram(mux_tree_tapbuf_size4_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_19_sram_inv[0:2]),
		.out(chany_bottom_out[22]));

	mux_tree_tapbuf_size4 mux_bottom_track_47 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[32], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size4_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_20_sram_inv[0:2]),
		.out(chany_bottom_out[23]));

	mux_tree_tapbuf_size4 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[33], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size4_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_21_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size4 mux_bottom_track_55 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[37], chanx_left_in[115]}),
		.sram(mux_tree_tapbuf_size4_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_22_sram_inv[0:2]),
		.out(chany_bottom_out[27]));

	mux_tree_tapbuf_size4 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[38], chanx_left_in[119]}),
		.sram(mux_tree_tapbuf_size4_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_23_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size4 mux_bottom_track_59 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[40], chanx_left_in[123]}),
		.sram(mux_tree_tapbuf_size4_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_24_sram_inv[0:2]),
		.out(chany_bottom_out[29]));

	mux_tree_tapbuf_size4 mux_bottom_track_61 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[41], chanx_left_in[127]}),
		.sram(mux_tree_tapbuf_size4_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_25_sram_inv[0:2]),
		.out(chany_bottom_out[30]));

	mux_tree_tapbuf_size4 mux_bottom_track_63 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[42], chanx_left_in[131]}),
		.sram(mux_tree_tapbuf_size4_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_26_sram_inv[0:2]),
		.out(chany_bottom_out[31]));

	mux_tree_tapbuf_size4 mux_bottom_track_65 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[44], chanx_left_in[135]}),
		.sram(mux_tree_tapbuf_size4_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_27_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size4 mux_bottom_track_67 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[45], chanx_left_in[139]}),
		.sram(mux_tree_tapbuf_size4_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_28_sram_inv[0:2]),
		.out(chany_bottom_out[33]));

	mux_tree_tapbuf_size4 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[49], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size4_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_29_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size4 mux_bottom_track_75 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[50], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size4_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_30_sram_inv[0:2]),
		.out(chany_bottom_out[37]));

	mux_tree_tapbuf_size4 mux_bottom_track_77 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[52], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size4_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_31_sram_inv[0:2]),
		.out(chany_bottom_out[38]));

	mux_tree_tapbuf_size4 mux_bottom_track_79 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[53], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size4_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_32_sram_inv[0:2]),
		.out(chany_bottom_out[39]));

	mux_tree_tapbuf_size4 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[54], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size4_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_33_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size4 mux_bottom_track_83 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[56], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size4_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_34_sram_inv[0:2]),
		.out(chany_bottom_out[41]));

	mux_tree_tapbuf_size4 mux_bottom_track_85 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[57], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size4_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_35_sram_inv[0:2]),
		.out(chany_bottom_out[42]));

	mux_tree_tapbuf_size4 mux_bottom_track_91 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[61], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size4_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_36_sram_inv[0:2]),
		.out(chany_bottom_out[45]));

	mux_tree_tapbuf_size4 mux_bottom_track_93 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[62], chanx_left_in[191]}),
		.sram(mux_tree_tapbuf_size4_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_37_sram_inv[0:2]),
		.out(chany_bottom_out[46]));

	mux_tree_tapbuf_size4 mux_bottom_track_95 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[64], chanx_left_in[195]}),
		.sram(mux_tree_tapbuf_size4_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_38_sram_inv[0:2]),
		.out(chany_bottom_out[47]));

	mux_tree_tapbuf_size4 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[65], chanx_left_in[199]}),
		.sram(mux_tree_tapbuf_size4_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_39_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size4 mux_bottom_track_99 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[66], chanx_left_in[203]}),
		.sram(mux_tree_tapbuf_size4_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_40_sram_inv[0:2]),
		.out(chany_bottom_out[49]));

	mux_tree_tapbuf_size4 mux_bottom_track_101 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[68], chanx_left_in[207]}),
		.sram(mux_tree_tapbuf_size4_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_41_sram_inv[0:2]),
		.out(chany_bottom_out[50]));

	mux_tree_tapbuf_size4 mux_bottom_track_103 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[69], chanx_left_in[211]}),
		.sram(mux_tree_tapbuf_size4_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_42_sram_inv[0:2]),
		.out(chany_bottom_out[51]));

	mux_tree_tapbuf_size4 mux_bottom_track_109 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[73], chanx_left_in[223]}),
		.sram(mux_tree_tapbuf_size4_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_43_sram_inv[0:2]),
		.out(chany_bottom_out[54]));

	mux_tree_tapbuf_size4 mux_bottom_track_111 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[74], chanx_left_in[227]}),
		.sram(mux_tree_tapbuf_size4_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_44_sram_inv[0:2]),
		.out(chany_bottom_out[55]));

	mux_tree_tapbuf_size4 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[76], chanx_left_in[231]}),
		.sram(mux_tree_tapbuf_size4_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_45_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size4 mux_bottom_track_115 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[77], chanx_left_in[235]}),
		.sram(mux_tree_tapbuf_size4_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_46_sram_inv[0:2]),
		.out(chany_bottom_out[57]));

	mux_tree_tapbuf_size4 mux_bottom_track_117 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[78], chanx_left_in[239]}),
		.sram(mux_tree_tapbuf_size4_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_47_sram_inv[0:2]),
		.out(chany_bottom_out[58]));

	mux_tree_tapbuf_size4 mux_bottom_track_119 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[80], chanx_left_in[243]}),
		.sram(mux_tree_tapbuf_size4_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_48_sram_inv[0:2]),
		.out(chany_bottom_out[59]));

	mux_tree_tapbuf_size4 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[81], chanx_left_in[247]}),
		.sram(mux_tree_tapbuf_size4_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_49_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size4 mux_bottom_track_127 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[85], chanx_left_in[259]}),
		.sram(mux_tree_tapbuf_size4_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_50_sram_inv[0:2]),
		.out(chany_bottom_out[63]));

	mux_tree_tapbuf_size4 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[86], chanx_left_in[263]}),
		.sram(mux_tree_tapbuf_size4_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_51_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size4 mux_bottom_track_131 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[88], chanx_left_in[267]}),
		.sram(mux_tree_tapbuf_size4_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_52_sram_inv[0:2]),
		.out(chany_bottom_out[65]));

	mux_tree_tapbuf_size4 mux_bottom_track_133 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[89], chanx_left_in[271]}),
		.sram(mux_tree_tapbuf_size4_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_53_sram_inv[0:2]),
		.out(chany_bottom_out[66]));

	mux_tree_tapbuf_size4 mux_bottom_track_135 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[90], chanx_left_in[275]}),
		.sram(mux_tree_tapbuf_size4_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_54_sram_inv[0:2]),
		.out(chany_bottom_out[67]));

	mux_tree_tapbuf_size4 mux_bottom_track_137 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[92], chanx_left_in[279]}),
		.sram(mux_tree_tapbuf_size4_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_55_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size4 mux_bottom_track_139 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[93], chanx_left_in[283]}),
		.sram(mux_tree_tapbuf_size4_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_56_sram_inv[0:2]),
		.out(chany_bottom_out[69]));

	mux_tree_tapbuf_size4 mux_bottom_track_145 (
		.in({chanx_right_in[281], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size4_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_57_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size4 mux_bottom_track_147 (
		.in({chanx_right_in[280], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size4_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_58_sram_inv[0:2]),
		.out(chany_bottom_out[73]));

	mux_tree_tapbuf_size4 mux_bottom_track_149 (
		.in({chanx_right_in[278], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size4_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_59_sram_inv[0:2]),
		.out(chany_bottom_out[74]));

	mux_tree_tapbuf_size4 mux_bottom_track_151 (
		.in({chanx_right_in[277], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size4_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_60_sram_inv[0:2]),
		.out(chany_bottom_out[75]));

	mux_tree_tapbuf_size4 mux_bottom_track_153 (
		.in({chanx_right_in[276], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size4_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_61_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size4 mux_bottom_track_155 (
		.in({chanx_right_in[274], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size4_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_62_sram_inv[0:2]),
		.out(chany_bottom_out[77]));

	mux_tree_tapbuf_size4 mux_bottom_track_157 (
		.in({chanx_right_in[273], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[105]}),
		.sram(mux_tree_tapbuf_size4_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_63_sram_inv[0:2]),
		.out(chany_bottom_out[78]));

	mux_tree_tapbuf_size4 mux_bottom_track_163 (
		.in({chanx_right_in[269], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[109]}),
		.sram(mux_tree_tapbuf_size4_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_64_sram_inv[0:2]),
		.out(chany_bottom_out[81]));

	mux_tree_tapbuf_size4 mux_bottom_track_165 (
		.in({chanx_right_in[268], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[110]}),
		.sram(mux_tree_tapbuf_size4_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_65_sram_inv[0:2]),
		.out(chany_bottom_out[82]));

	mux_tree_tapbuf_size4 mux_bottom_track_167 (
		.in({chanx_right_in[266], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[112]}),
		.sram(mux_tree_tapbuf_size4_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_66_sram_inv[0:2]),
		.out(chany_bottom_out[83]));

	mux_tree_tapbuf_size4 mux_bottom_track_169 (
		.in({chanx_right_in[265], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[113]}),
		.sram(mux_tree_tapbuf_size4_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_67_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size4 mux_bottom_track_171 (
		.in({chanx_right_in[264], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[114]}),
		.sram(mux_tree_tapbuf_size4_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_68_sram_inv[0:2]),
		.out(chany_bottom_out[85]));

	mux_tree_tapbuf_size4 mux_bottom_track_173 (
		.in({chanx_right_in[262], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[116]}),
		.sram(mux_tree_tapbuf_size4_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_69_sram_inv[0:2]),
		.out(chany_bottom_out[86]));

	mux_tree_tapbuf_size4 mux_bottom_track_175 (
		.in({chanx_right_in[261], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[117]}),
		.sram(mux_tree_tapbuf_size4_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_70_sram_inv[0:2]),
		.out(chany_bottom_out[87]));

	mux_tree_tapbuf_size4 mux_bottom_track_181 (
		.in({chanx_right_in[257], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[121]}),
		.sram(mux_tree_tapbuf_size4_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_71_sram_inv[0:2]),
		.out(chany_bottom_out[90]));

	mux_tree_tapbuf_size4 mux_bottom_track_183 (
		.in({chanx_right_in[256], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[122]}),
		.sram(mux_tree_tapbuf_size4_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_72_sram_inv[0:2]),
		.out(chany_bottom_out[91]));

	mux_tree_tapbuf_size4 mux_bottom_track_185 (
		.in({chanx_right_in[254], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[124]}),
		.sram(mux_tree_tapbuf_size4_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_73_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size4 mux_bottom_track_187 (
		.in({chanx_right_in[253], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[125]}),
		.sram(mux_tree_tapbuf_size4_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_74_sram_inv[0:2]),
		.out(chany_bottom_out[93]));

	mux_tree_tapbuf_size4 mux_bottom_track_189 (
		.in({chanx_right_in[252], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[126]}),
		.sram(mux_tree_tapbuf_size4_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_75_sram_inv[0:2]),
		.out(chany_bottom_out[94]));

	mux_tree_tapbuf_size4 mux_bottom_track_191 (
		.in({chanx_right_in[250], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size4_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_76_sram_inv[0:2]),
		.out(chany_bottom_out[95]));

	mux_tree_tapbuf_size4 mux_bottom_track_193 (
		.in({chanx_right_in[249], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size4_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_77_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size4 mux_bottom_track_199 (
		.in({chanx_right_in[245], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size4_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_78_sram_inv[0:2]),
		.out(chany_bottom_out[99]));

	mux_tree_tapbuf_size4 mux_bottom_track_201 (
		.in({chanx_right_in[244], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size4_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_79_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size4 mux_bottom_track_203 (
		.in({chanx_right_in[242], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size4_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_80_sram_inv[0:2]),
		.out(chany_bottom_out[101]));

	mux_tree_tapbuf_size4 mux_bottom_track_205 (
		.in({chanx_right_in[241], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size4_81_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_81_sram_inv[0:2]),
		.out(chany_bottom_out[102]));

	mux_tree_tapbuf_size4 mux_bottom_track_207 (
		.in({chanx_right_in[240], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size4_82_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_82_sram_inv[0:2]),
		.out(chany_bottom_out[103]));

	mux_tree_tapbuf_size4 mux_bottom_track_209 (
		.in({chanx_right_in[238], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size4_83_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_83_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size4 mux_bottom_track_211 (
		.in({chanx_right_in[237], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size4_84_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_84_sram_inv[0:2]),
		.out(chany_bottom_out[105]));

	mux_tree_tapbuf_size4 mux_bottom_track_217 (
		.in({chanx_right_in[233], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size4_85_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_85_sram_inv[0:2]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size4 mux_bottom_track_219 (
		.in({chanx_right_in[232], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size4_86_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_86_sram_inv[0:2]),
		.out(chany_bottom_out[109]));

	mux_tree_tapbuf_size4 mux_bottom_track_221 (
		.in({chanx_right_in[230], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size4_87_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_87_sram_inv[0:2]),
		.out(chany_bottom_out[110]));

	mux_tree_tapbuf_size4 mux_bottom_track_223 (
		.in({chanx_right_in[229], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size4_88_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_88_sram_inv[0:2]),
		.out(chany_bottom_out[111]));

	mux_tree_tapbuf_size4 mux_bottom_track_225 (
		.in({chanx_right_in[228], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size4_89_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_89_sram_inv[0:2]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size4 mux_bottom_track_227 (
		.in({chanx_right_in[226], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size4_90_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_90_sram_inv[0:2]),
		.out(chany_bottom_out[113]));

	mux_tree_tapbuf_size4 mux_bottom_track_229 (
		.in({chanx_right_in[225], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size4_91_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_91_sram_inv[0:2]),
		.out(chany_bottom_out[114]));

	mux_tree_tapbuf_size4 mux_bottom_track_235 (
		.in({chanx_right_in[221], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size4_92_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_92_sram_inv[0:2]),
		.out(chany_bottom_out[117]));

	mux_tree_tapbuf_size4 mux_bottom_track_237 (
		.in({chanx_right_in[220], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size4_93_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_93_sram_inv[0:2]),
		.out(chany_bottom_out[118]));

	mux_tree_tapbuf_size4 mux_bottom_track_239 (
		.in({chanx_right_in[218], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size4_94_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_94_sram_inv[0:2]),
		.out(chany_bottom_out[119]));

	mux_tree_tapbuf_size4 mux_bottom_track_241 (
		.in({chanx_right_in[217], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size4_95_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_95_sram_inv[0:2]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size4 mux_bottom_track_243 (
		.in({chanx_right_in[216], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size4_96_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_96_sram_inv[0:2]),
		.out(chany_bottom_out[121]));

	mux_tree_tapbuf_size4 mux_bottom_track_245 (
		.in({chanx_right_in[214], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size4_97_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_97_sram_inv[0:2]),
		.out(chany_bottom_out[122]));

	mux_tree_tapbuf_size4 mux_bottom_track_247 (
		.in({chanx_right_in[213], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size4_98_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_98_sram_inv[0:2]),
		.out(chany_bottom_out[123]));

	mux_tree_tapbuf_size4 mux_bottom_track_253 (
		.in({chanx_right_in[209], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size4_99_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_99_sram_inv[0:2]),
		.out(chany_bottom_out[126]));

	mux_tree_tapbuf_size4 mux_bottom_track_255 (
		.in({chanx_right_in[208], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size4_100_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_100_sram_inv[0:2]),
		.out(chany_bottom_out[127]));

	mux_tree_tapbuf_size4 mux_bottom_track_257 (
		.in({chanx_right_in[206], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size4_101_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_101_sram_inv[0:2]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size4 mux_bottom_track_259 (
		.in({chanx_right_in[205], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size4_102_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_102_sram_inv[0:2]),
		.out(chany_bottom_out[129]));

	mux_tree_tapbuf_size4 mux_bottom_track_261 (
		.in({chanx_right_in[204], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size4_103_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_103_sram_inv[0:2]),
		.out(chany_bottom_out[130]));

	mux_tree_tapbuf_size4 mux_bottom_track_263 (
		.in({chanx_right_in[202], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size4_104_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_104_sram_inv[0:2]),
		.out(chany_bottom_out[131]));

	mux_tree_tapbuf_size4 mux_bottom_track_265 (
		.in({chanx_right_in[201], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size4_105_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_105_sram_inv[0:2]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size4 mux_bottom_track_271 (
		.in({chanx_right_in[197], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size4_106_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_106_sram_inv[0:2]),
		.out(chany_bottom_out[135]));

	mux_tree_tapbuf_size4 mux_bottom_track_273 (
		.in({chanx_right_in[196], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size4_107_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_107_sram_inv[0:2]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size4 mux_bottom_track_275 (
		.in({chanx_right_in[194], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size4_108_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_108_sram_inv[0:2]),
		.out(chany_bottom_out[137]));

	mux_tree_tapbuf_size4 mux_bottom_track_277 (
		.in({chanx_right_in[193], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size4_109_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_109_sram_inv[0:2]),
		.out(chany_bottom_out[138]));

	mux_tree_tapbuf_size4 mux_bottom_track_279 (
		.in({chanx_right_in[192], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size4_110_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_110_sram_inv[0:2]),
		.out(chany_bottom_out[139]));

	mux_tree_tapbuf_size4 mux_bottom_track_281 (
		.in({chanx_right_in[190], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size4_111_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_111_sram_inv[0:2]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size4 mux_bottom_track_283 (
		.in({chanx_right_in[189], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[189]}),
		.sram(mux_tree_tapbuf_size4_112_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_112_sram_inv[0:2]),
		.out(chany_bottom_out[141]));

	mux_tree_tapbuf_size4 mux_bottom_track_289 (
		.in({chanx_right_in[185], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[193]}),
		.sram(mux_tree_tapbuf_size4_113_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_113_sram_inv[0:2]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size4 mux_bottom_track_291 (
		.in({chanx_right_in[184], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[194]}),
		.sram(mux_tree_tapbuf_size4_114_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_114_sram_inv[0:2]),
		.out(chany_bottom_out[145]));

	mux_tree_tapbuf_size4 mux_bottom_track_293 (
		.in({chanx_right_in[182], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[196]}),
		.sram(mux_tree_tapbuf_size4_115_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_115_sram_inv[0:2]),
		.out(chany_bottom_out[146]));

	mux_tree_tapbuf_size4 mux_bottom_track_295 (
		.in({chanx_right_in[181], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[197]}),
		.sram(mux_tree_tapbuf_size4_116_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_116_sram_inv[0:2]),
		.out(chany_bottom_out[147]));

	mux_tree_tapbuf_size4 mux_bottom_track_297 (
		.in({chanx_right_in[180], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[198]}),
		.sram(mux_tree_tapbuf_size4_117_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_117_sram_inv[0:2]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size4 mux_bottom_track_299 (
		.in({chanx_right_in[178], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[200]}),
		.sram(mux_tree_tapbuf_size4_118_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_118_sram_inv[0:2]),
		.out(chany_bottom_out[149]));

	mux_tree_tapbuf_size4 mux_bottom_track_301 (
		.in({chanx_right_in[177], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[201]}),
		.sram(mux_tree_tapbuf_size4_119_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_119_sram_inv[0:2]),
		.out(chany_bottom_out[150]));

	mux_tree_tapbuf_size4 mux_bottom_track_307 (
		.in({chanx_right_in[173], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[205]}),
		.sram(mux_tree_tapbuf_size4_120_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_120_sram_inv[0:2]),
		.out(chany_bottom_out[153]));

	mux_tree_tapbuf_size4 mux_bottom_track_309 (
		.in({chanx_right_in[172], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[206]}),
		.sram(mux_tree_tapbuf_size4_121_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_121_sram_inv[0:2]),
		.out(chany_bottom_out[154]));

	mux_tree_tapbuf_size4 mux_bottom_track_311 (
		.in({chanx_right_in[170], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[208]}),
		.sram(mux_tree_tapbuf_size4_122_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_122_sram_inv[0:2]),
		.out(chany_bottom_out[155]));

	mux_tree_tapbuf_size4 mux_bottom_track_313 (
		.in({chanx_right_in[169], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[209]}),
		.sram(mux_tree_tapbuf_size4_123_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_123_sram_inv[0:2]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size4 mux_bottom_track_315 (
		.in({chanx_right_in[168], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[210]}),
		.sram(mux_tree_tapbuf_size4_124_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_124_sram_inv[0:2]),
		.out(chany_bottom_out[157]));

	mux_tree_tapbuf_size4 mux_bottom_track_317 (
		.in({chanx_right_in[166], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[212]}),
		.sram(mux_tree_tapbuf_size4_125_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_125_sram_inv[0:2]),
		.out(chany_bottom_out[158]));

	mux_tree_tapbuf_size4 mux_bottom_track_319 (
		.in({chanx_right_in[165], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[213]}),
		.sram(mux_tree_tapbuf_size4_126_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_126_sram_inv[0:2]),
		.out(chany_bottom_out[159]));

	mux_tree_tapbuf_size4 mux_bottom_track_325 (
		.in({chanx_right_in[161], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[217]}),
		.sram(mux_tree_tapbuf_size4_127_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_127_sram_inv[0:2]),
		.out(chany_bottom_out[162]));

	mux_tree_tapbuf_size4 mux_bottom_track_327 (
		.in({chanx_right_in[160], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[218]}),
		.sram(mux_tree_tapbuf_size4_128_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_128_sram_inv[0:2]),
		.out(chany_bottom_out[163]));

	mux_tree_tapbuf_size4 mux_bottom_track_329 (
		.in({chanx_right_in[158], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[220]}),
		.sram(mux_tree_tapbuf_size4_129_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_129_sram_inv[0:2]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size4 mux_bottom_track_331 (
		.in({chanx_right_in[157], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[221]}),
		.sram(mux_tree_tapbuf_size4_130_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_130_sram_inv[0:2]),
		.out(chany_bottom_out[165]));

	mux_tree_tapbuf_size4 mux_bottom_track_333 (
		.in({chanx_right_in[156], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[222]}),
		.sram(mux_tree_tapbuf_size4_131_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_131_sram_inv[0:2]),
		.out(chany_bottom_out[166]));

	mux_tree_tapbuf_size4 mux_bottom_track_335 (
		.in({chanx_right_in[154], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[224]}),
		.sram(mux_tree_tapbuf_size4_132_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_132_sram_inv[0:2]),
		.out(chany_bottom_out[167]));

	mux_tree_tapbuf_size4 mux_bottom_track_337 (
		.in({chanx_right_in[153], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[225]}),
		.sram(mux_tree_tapbuf_size4_133_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_133_sram_inv[0:2]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size4 mux_bottom_track_343 (
		.in({chanx_right_in[149], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[229]}),
		.sram(mux_tree_tapbuf_size4_134_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_134_sram_inv[0:2]),
		.out(chany_bottom_out[171]));

	mux_tree_tapbuf_size4 mux_bottom_track_345 (
		.in({chanx_right_in[148], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[230]}),
		.sram(mux_tree_tapbuf_size4_135_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_135_sram_inv[0:2]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size4 mux_bottom_track_347 (
		.in({chanx_right_in[146], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[232]}),
		.sram(mux_tree_tapbuf_size4_136_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_136_sram_inv[0:2]),
		.out(chany_bottom_out[173]));

	mux_tree_tapbuf_size4 mux_bottom_track_349 (
		.in({chanx_right_in[145], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[233]}),
		.sram(mux_tree_tapbuf_size4_137_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_137_sram_inv[0:2]),
		.out(chany_bottom_out[174]));

	mux_tree_tapbuf_size4 mux_bottom_track_351 (
		.in({chanx_right_in[144], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[234]}),
		.sram(mux_tree_tapbuf_size4_138_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_138_sram_inv[0:2]),
		.out(chany_bottom_out[175]));

	mux_tree_tapbuf_size4 mux_bottom_track_353 (
		.in({chanx_right_in[142], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[236]}),
		.sram(mux_tree_tapbuf_size4_139_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_139_sram_inv[0:2]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size4 mux_bottom_track_355 (
		.in({chanx_right_in[141], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[237]}),
		.sram(mux_tree_tapbuf_size4_140_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_140_sram_inv[0:2]),
		.out(chany_bottom_out[177]));

	mux_tree_tapbuf_size4 mux_bottom_track_361 (
		.in({chanx_right_in[137], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[241]}),
		.sram(mux_tree_tapbuf_size4_141_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_141_sram_inv[0:2]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size4 mux_bottom_track_363 (
		.in({chanx_right_in[136], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[242]}),
		.sram(mux_tree_tapbuf_size4_142_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_142_sram_inv[0:2]),
		.out(chany_bottom_out[181]));

	mux_tree_tapbuf_size4 mux_bottom_track_365 (
		.in({chanx_right_in[134], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[244]}),
		.sram(mux_tree_tapbuf_size4_143_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_143_sram_inv[0:2]),
		.out(chany_bottom_out[182]));

	mux_tree_tapbuf_size4 mux_bottom_track_367 (
		.in({chanx_right_in[133], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[245]}),
		.sram(mux_tree_tapbuf_size4_144_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_144_sram_inv[0:2]),
		.out(chany_bottom_out[183]));

	mux_tree_tapbuf_size4 mux_bottom_track_369 (
		.in({chanx_right_in[132], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[246]}),
		.sram(mux_tree_tapbuf_size4_145_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_145_sram_inv[0:2]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size4 mux_bottom_track_371 (
		.in({chanx_right_in[130], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[248]}),
		.sram(mux_tree_tapbuf_size4_146_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_146_sram_inv[0:2]),
		.out(chany_bottom_out[185]));

	mux_tree_tapbuf_size4 mux_bottom_track_373 (
		.in({chanx_right_in[129], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[249]}),
		.sram(mux_tree_tapbuf_size4_147_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_147_sram_inv[0:2]),
		.out(chany_bottom_out[186]));

	mux_tree_tapbuf_size4 mux_bottom_track_379 (
		.in({chanx_right_in[125], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[253]}),
		.sram(mux_tree_tapbuf_size4_148_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_148_sram_inv[0:2]),
		.out(chany_bottom_out[189]));

	mux_tree_tapbuf_size4 mux_bottom_track_381 (
		.in({chanx_right_in[124], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[254]}),
		.sram(mux_tree_tapbuf_size4_149_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_149_sram_inv[0:2]),
		.out(chany_bottom_out[190]));

	mux_tree_tapbuf_size4 mux_bottom_track_383 (
		.in({chanx_right_in[122], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[256]}),
		.sram(mux_tree_tapbuf_size4_150_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_150_sram_inv[0:2]),
		.out(chany_bottom_out[191]));

	mux_tree_tapbuf_size4 mux_bottom_track_385 (
		.in({chanx_right_in[121], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[257]}),
		.sram(mux_tree_tapbuf_size4_151_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_151_sram_inv[0:2]),
		.out(chany_bottom_out[192]));

	mux_tree_tapbuf_size4 mux_bottom_track_387 (
		.in({chanx_right_in[120], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[258]}),
		.sram(mux_tree_tapbuf_size4_152_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_152_sram_inv[0:2]),
		.out(chany_bottom_out[193]));

	mux_tree_tapbuf_size4 mux_bottom_track_389 (
		.in({chanx_right_in[118], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[260]}),
		.sram(mux_tree_tapbuf_size4_153_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_153_sram_inv[0:2]),
		.out(chany_bottom_out[194]));

	mux_tree_tapbuf_size4 mux_bottom_track_391 (
		.in({chanx_right_in[117], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[261]}),
		.sram(mux_tree_tapbuf_size4_154_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_154_sram_inv[0:2]),
		.out(chany_bottom_out[195]));

	mux_tree_tapbuf_size4 mux_bottom_track_397 (
		.in({chanx_right_in[113], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[265]}),
		.sram(mux_tree_tapbuf_size4_155_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_155_sram_inv[0:2]),
		.out(chany_bottom_out[198]));

	mux_tree_tapbuf_size4 mux_bottom_track_399 (
		.in({chanx_right_in[112], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[266]}),
		.sram(mux_tree_tapbuf_size4_156_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_156_sram_inv[0:2]),
		.out(chany_bottom_out[199]));

	mux_tree_tapbuf_size4 mux_bottom_track_401 (
		.in({chanx_right_in[110], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[268]}),
		.sram(mux_tree_tapbuf_size4_157_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_157_sram_inv[0:2]),
		.out(chany_bottom_out[200]));

	mux_tree_tapbuf_size4 mux_bottom_track_403 (
		.in({chanx_right_in[109], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[269]}),
		.sram(mux_tree_tapbuf_size4_158_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_158_sram_inv[0:2]),
		.out(chany_bottom_out[201]));

	mux_tree_tapbuf_size4 mux_bottom_track_405 (
		.in({chanx_right_in[108], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[270]}),
		.sram(mux_tree_tapbuf_size4_159_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_159_sram_inv[0:2]),
		.out(chany_bottom_out[202]));

	mux_tree_tapbuf_size4 mux_bottom_track_407 (
		.in({chanx_right_in[106], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[272]}),
		.sram(mux_tree_tapbuf_size4_160_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_160_sram_inv[0:2]),
		.out(chany_bottom_out[203]));

	mux_tree_tapbuf_size4 mux_bottom_track_409 (
		.in({chanx_right_in[105], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[273]}),
		.sram(mux_tree_tapbuf_size4_161_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_161_sram_inv[0:2]),
		.out(chany_bottom_out[204]));

	mux_tree_tapbuf_size4 mux_bottom_track_415 (
		.in({chanx_right_in[101], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[277]}),
		.sram(mux_tree_tapbuf_size4_162_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_162_sram_inv[0:2]),
		.out(chany_bottom_out[207]));

	mux_tree_tapbuf_size4 mux_bottom_track_417 (
		.in({chanx_right_in[100], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[278]}),
		.sram(mux_tree_tapbuf_size4_163_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_163_sram_inv[0:2]),
		.out(chany_bottom_out[208]));

	mux_tree_tapbuf_size4 mux_bottom_track_419 (
		.in({chanx_right_in[98], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[280]}),
		.sram(mux_tree_tapbuf_size4_164_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_164_sram_inv[0:2]),
		.out(chany_bottom_out[209]));

	mux_tree_tapbuf_size4 mux_bottom_track_421 (
		.in({chanx_right_in[97], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[281]}),
		.sram(mux_tree_tapbuf_size4_165_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_165_sram_inv[0:2]),
		.out(chany_bottom_out[210]));

	mux_tree_tapbuf_size4 mux_bottom_track_423 (
		.in({chanx_right_in[96], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[282]}),
		.sram(mux_tree_tapbuf_size4_166_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_166_sram_inv[0:2]),
		.out(chany_bottom_out[211]));

	mux_tree_tapbuf_size4 mux_bottom_track_425 (
		.in({chanx_right_in[94], chanx_right_in[284], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_167_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_167_sram_inv[0:2]),
		.out(chany_bottom_out[212]));

	mux_tree_tapbuf_size4 mux_bottom_track_427 (
		.in({chanx_right_in[93], chanx_right_in[283], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_168_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_168_sram_inv[0:2]),
		.out(chany_bottom_out[213]));

	mux_tree_tapbuf_size4 mux_bottom_track_433 (
		.in({chanx_right_in[89], chanx_right_in[271], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_169_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_169_sram_inv[0:2]),
		.out(chany_bottom_out[216]));

	mux_tree_tapbuf_size4 mux_bottom_track_435 (
		.in({chanx_right_in[88], chanx_right_in[267], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_170_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_170_sram_inv[0:2]),
		.out(chany_bottom_out[217]));

	mux_tree_tapbuf_size4 mux_bottom_track_437 (
		.in({chanx_right_in[86], chanx_right_in[263], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_171_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_171_sram_inv[0:2]),
		.out(chany_bottom_out[218]));

	mux_tree_tapbuf_size4 mux_bottom_track_439 (
		.in({chanx_right_in[85], chanx_right_in[259], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_172_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_172_sram_inv[0:2]),
		.out(chany_bottom_out[219]));

	mux_tree_tapbuf_size4 mux_bottom_track_441 (
		.in({chanx_right_in[84], chanx_right_in[255], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_173_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_173_sram_inv[0:2]),
		.out(chany_bottom_out[220]));

	mux_tree_tapbuf_size4 mux_bottom_track_443 (
		.in({chanx_right_in[82], chanx_right_in[251], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_174_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_174_sram_inv[0:2]),
		.out(chany_bottom_out[221]));

	mux_tree_tapbuf_size4 mux_bottom_track_445 (
		.in({chanx_right_in[81], chanx_right_in[247], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_175_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_175_sram_inv[0:2]),
		.out(chany_bottom_out[222]));

	mux_tree_tapbuf_size4 mux_bottom_track_451 (
		.in({chanx_right_in[77], chanx_right_in[235], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_176_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_176_sram_inv[0:2]),
		.out(chany_bottom_out[225]));

	mux_tree_tapbuf_size4 mux_bottom_track_453 (
		.in({chanx_right_in[76], chanx_right_in[231], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_177_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_177_sram_inv[0:2]),
		.out(chany_bottom_out[226]));

	mux_tree_tapbuf_size4 mux_bottom_track_455 (
		.in({chanx_right_in[74], chanx_right_in[227], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_178_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_178_sram_inv[0:2]),
		.out(chany_bottom_out[227]));

	mux_tree_tapbuf_size4 mux_bottom_track_457 (
		.in({chanx_right_in[73], chanx_right_in[223], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_179_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_179_sram_inv[0:2]),
		.out(chany_bottom_out[228]));

	mux_tree_tapbuf_size4 mux_bottom_track_459 (
		.in({chanx_right_in[72], chanx_right_in[219], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_180_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_180_sram_inv[0:2]),
		.out(chany_bottom_out[229]));

	mux_tree_tapbuf_size4 mux_bottom_track_461 (
		.in({chanx_right_in[70], chanx_right_in[215], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_181_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_181_sram_inv[0:2]),
		.out(chany_bottom_out[230]));

	mux_tree_tapbuf_size4 mux_bottom_track_463 (
		.in({chanx_right_in[69], chanx_right_in[211], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_182_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_182_sram_inv[0:2]),
		.out(chany_bottom_out[231]));

	mux_tree_tapbuf_size4 mux_bottom_track_469 (
		.in({chanx_right_in[65], chanx_right_in[199], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_183_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_183_sram_inv[0:2]),
		.out(chany_bottom_out[234]));

	mux_tree_tapbuf_size4 mux_bottom_track_471 (
		.in({chanx_right_in[64], chanx_right_in[195], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_184_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_184_sram_inv[0:2]),
		.out(chany_bottom_out[235]));

	mux_tree_tapbuf_size4 mux_bottom_track_473 (
		.in({chanx_right_in[62], chanx_right_in[191], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_185_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_185_sram_inv[0:2]),
		.out(chany_bottom_out[236]));

	mux_tree_tapbuf_size4 mux_bottom_track_475 (
		.in({chanx_right_in[61], chanx_right_in[187], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_186_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_186_sram_inv[0:2]),
		.out(chany_bottom_out[237]));

	mux_tree_tapbuf_size4 mux_bottom_track_477 (
		.in({chanx_right_in[60], chanx_right_in[183], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_187_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_187_sram_inv[0:2]),
		.out(chany_bottom_out[238]));

	mux_tree_tapbuf_size4 mux_bottom_track_479 (
		.in({chanx_right_in[58], chanx_right_in[179], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_188_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_188_sram_inv[0:2]),
		.out(chany_bottom_out[239]));

	mux_tree_tapbuf_size4 mux_bottom_track_481 (
		.in({chanx_right_in[57], chanx_right_in[175], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_189_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_189_sram_inv[0:2]),
		.out(chany_bottom_out[240]));

	mux_tree_tapbuf_size4 mux_bottom_track_487 (
		.in({chanx_right_in[53], chanx_right_in[163], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_190_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_190_sram_inv[0:2]),
		.out(chany_bottom_out[243]));

	mux_tree_tapbuf_size4 mux_bottom_track_489 (
		.in({chanx_right_in[52], chanx_right_in[159], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_191_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_191_sram_inv[0:2]),
		.out(chany_bottom_out[244]));

	mux_tree_tapbuf_size4 mux_bottom_track_491 (
		.in({chanx_right_in[50], chanx_right_in[155], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_192_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_192_sram_inv[0:2]),
		.out(chany_bottom_out[245]));

	mux_tree_tapbuf_size4 mux_bottom_track_493 (
		.in({chanx_right_in[49], chanx_right_in[151], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_193_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_193_sram_inv[0:2]),
		.out(chany_bottom_out[246]));

	mux_tree_tapbuf_size4 mux_bottom_track_495 (
		.in({chanx_right_in[48], chanx_right_in[147], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_194_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_194_sram_inv[0:2]),
		.out(chany_bottom_out[247]));

	mux_tree_tapbuf_size4 mux_bottom_track_497 (
		.in({chanx_right_in[46], chanx_right_in[143], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_195_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_195_sram_inv[0:2]),
		.out(chany_bottom_out[248]));

	mux_tree_tapbuf_size4 mux_bottom_track_499 (
		.in({chanx_right_in[45], chanx_right_in[139], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_196_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_196_sram_inv[0:2]),
		.out(chany_bottom_out[249]));

	mux_tree_tapbuf_size4 mux_bottom_track_505 (
		.in({chanx_right_in[41], chanx_right_in[127], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_197_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_197_sram_inv[0:2]),
		.out(chany_bottom_out[252]));

	mux_tree_tapbuf_size4 mux_bottom_track_507 (
		.in({chanx_right_in[40], chanx_right_in[123], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_198_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_198_sram_inv[0:2]),
		.out(chany_bottom_out[253]));

	mux_tree_tapbuf_size4 mux_bottom_track_509 (
		.in({chanx_right_in[38], chanx_right_in[119], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_199_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_199_sram_inv[0:2]),
		.out(chany_bottom_out[254]));

	mux_tree_tapbuf_size4 mux_bottom_track_511 (
		.in({chanx_right_in[37], chanx_right_in[115], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_200_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_200_sram_inv[0:2]),
		.out(chany_bottom_out[255]));

	mux_tree_tapbuf_size4 mux_bottom_track_513 (
		.in({chanx_right_in[36], chanx_right_in[111], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_201_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_201_sram_inv[0:2]),
		.out(chany_bottom_out[256]));

	mux_tree_tapbuf_size4 mux_bottom_track_515 (
		.in({chanx_right_in[34], chanx_right_in[107], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_202_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_202_sram_inv[0:2]),
		.out(chany_bottom_out[257]));

	mux_tree_tapbuf_size4 mux_bottom_track_517 (
		.in({chanx_right_in[33], chanx_right_in[103], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_203_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_203_sram_inv[0:2]),
		.out(chany_bottom_out[258]));

	mux_tree_tapbuf_size4 mux_bottom_track_523 (
		.in({chanx_right_in[29], chanx_right_in[91], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_204_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_204_sram_inv[0:2]),
		.out(chany_bottom_out[261]));

	mux_tree_tapbuf_size4 mux_bottom_track_525 (
		.in({chanx_right_in[28], chanx_right_in[87], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_205_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_205_sram_inv[0:2]),
		.out(chany_bottom_out[262]));

	mux_tree_tapbuf_size4 mux_bottom_track_527 (
		.in({chanx_right_in[26], chanx_right_in[83], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_206_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_206_sram_inv[0:2]),
		.out(chany_bottom_out[263]));

	mux_tree_tapbuf_size4 mux_bottom_track_529 (
		.in({chanx_right_in[25], chanx_right_in[79], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_207_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_207_sram_inv[0:2]),
		.out(chany_bottom_out[264]));

	mux_tree_tapbuf_size4 mux_bottom_track_531 (
		.in({chanx_right_in[24], chanx_right_in[75], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_208_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_208_sram_inv[0:2]),
		.out(chany_bottom_out[265]));

	mux_tree_tapbuf_size4 mux_bottom_track_533 (
		.in({chanx_right_in[22], chanx_right_in[71], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_209_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_209_sram_inv[0:2]),
		.out(chany_bottom_out[266]));

	mux_tree_tapbuf_size4 mux_bottom_track_535 (
		.in({chanx_right_in[21], chanx_right_in[67], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_210_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_210_sram_inv[0:2]),
		.out(chany_bottom_out[267]));

	mux_tree_tapbuf_size4 mux_bottom_track_541 (
		.in({chanx_right_in[17], chanx_right_in[55], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_211_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_211_sram_inv[0:2]),
		.out(chany_bottom_out[270]));

	mux_tree_tapbuf_size4 mux_bottom_track_543 (
		.in({chanx_right_in[16], chanx_right_in[51], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_212_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_212_sram_inv[0:2]),
		.out(chany_bottom_out[271]));

	mux_tree_tapbuf_size4 mux_bottom_track_545 (
		.in({chanx_right_in[14], chanx_right_in[47], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_213_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_213_sram_inv[0:2]),
		.out(chany_bottom_out[272]));

	mux_tree_tapbuf_size4 mux_bottom_track_547 (
		.in({chanx_right_in[13], chanx_right_in[43], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_214_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_214_sram_inv[0:2]),
		.out(chany_bottom_out[273]));

	mux_tree_tapbuf_size4 mux_bottom_track_549 (
		.in({chanx_right_in[12], chanx_right_in[39], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_215_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_215_sram_inv[0:2]),
		.out(chany_bottom_out[274]));

	mux_tree_tapbuf_size4 mux_bottom_track_551 (
		.in({chanx_right_in[10], chanx_right_in[35], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_216_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_216_sram_inv[0:2]),
		.out(chany_bottom_out[275]));

	mux_tree_tapbuf_size4 mux_bottom_track_553 (
		.in({chanx_right_in[9], chanx_right_in[31], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_217_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_217_sram_inv[0:2]),
		.out(chany_bottom_out[276]));

	mux_tree_tapbuf_size4 mux_bottom_track_559 (
		.in({chanx_right_in[5], chanx_right_in[19], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_218_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_218_sram_inv[0:2]),
		.out(chany_bottom_out[279]));

	mux_tree_tapbuf_size4 mux_bottom_track_561 (
		.in({chanx_right_in[4], chanx_right_in[15], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_219_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_219_sram_inv[0:2]),
		.out(chany_bottom_out[280]));

	mux_tree_tapbuf_size4 mux_bottom_track_563 (
		.in({chanx_right_in[2], chanx_right_in[11], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_220_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_220_sram_inv[0:2]),
		.out(chany_bottom_out[281]));

	mux_tree_tapbuf_size4 mux_bottom_track_565 (
		.in({chanx_right_in[1], chanx_right_in[7], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_221_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_221_sram_inv[0:2]),
		.out(chany_bottom_out[282]));

	mux_tree_tapbuf_size4 mux_bottom_track_567 (
		.in({chanx_right_in[0], chanx_right_in[3], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_222_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_222_sram_inv[0:2]),
		.out(chany_bottom_out[283]));

	mux_tree_tapbuf_size4 mux_bottom_track_569 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[0], chanx_left_in[3]}),
		.sram(mux_tree_tapbuf_size4_223_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_223_sram_inv[0:2]),
		.out(chany_bottom_out[284]));

	mux_tree_tapbuf_size4 mux_left_track_561 (
		.in({chany_bottom_in[69], chany_bottom_in[141], chany_bottom_in[213], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_224_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_224_sram_inv[0:2]),
		.out(chanx_left_out[280]));

	mux_tree_tapbuf_size4 mux_left_track_569 (
		.in({chany_bottom_in[70], chany_bottom_in[142], chany_bottom_in[214], left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_225_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_225_sram_inv[0:2]),
		.out(chanx_left_out[284]));

	mux_tree_tapbuf_size4_mem mem_right_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_7_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_8_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_9_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_10_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_11_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_12_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_13_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_14_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_15_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_16_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_17_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_18_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_19_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_20_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_21_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_22_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_23_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_24_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_25_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_26_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_27_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_28_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_29_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_30_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_31_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_32_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_33_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_34_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_35_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_36_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_37_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_38_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_39_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_40_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_41_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_42_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_43_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_44_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_45_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_46_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_47_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_48_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_49_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_50_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_51_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_52_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_53_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_54_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_55_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_56_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_57_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_58_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_59_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_60_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_61_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_62_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_63_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_64_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_65_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_66_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_67_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_68_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_69_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_70_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_71_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_72_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_73_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_74_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_75_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_76_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_77_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_78_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_79_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_80_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_81_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_81_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_82_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_82_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_83_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_83_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_84_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_84_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_85_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_85_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_219 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_86_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_86_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_221 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_87_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_87_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_223 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_88_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_88_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_89_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_89_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_227 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_90_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_90_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_229 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_91_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_91_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_235 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_92_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_92_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_237 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_93_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_93_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_239 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_94_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_94_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_95_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_95_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_243 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_96_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_96_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_245 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_97_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_97_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_247 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_98_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_98_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_253 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_99_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_99_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_255 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_100_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_100_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_101_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_101_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_259 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_102_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_102_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_261 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_103_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_103_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_263 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_104_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_104_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_105_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_105_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_271 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_106_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_106_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_107_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_107_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_275 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_108_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_108_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_277 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_109_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_109_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_279 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_110_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_110_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_111_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_111_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_283 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_112_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_112_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_113_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_113_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_291 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_114_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_114_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_293 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_115_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_115_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_295 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_116_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_116_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_117_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_117_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_299 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_118_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_118_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_301 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_119_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_119_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_307 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_120_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_120_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_309 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_121_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_121_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_311 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_122_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_122_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_123_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_123_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_315 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_124_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_124_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_317 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_125_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_125_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_319 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_126_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_126_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_325 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_127_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_127_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_327 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_128_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_128_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_129_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_129_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_331 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_130_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_130_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_333 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_131_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_131_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_335 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_132_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_132_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_133_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_133_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_343 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_134_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_134_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_135_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_135_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_347 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_136_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_136_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_349 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_137_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_137_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_351 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_138_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_138_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_139_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_139_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_355 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_140_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_140_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_141_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_141_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_363 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_142_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_142_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_365 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_143_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_143_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_367 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_144_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_144_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_145_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_145_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_371 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_146_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_146_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_373 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_147_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_147_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_379 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_148_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_148_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_381 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_149_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_149_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_383 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_150_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_150_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_151_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_151_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_387 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_152_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_152_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_389 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_153_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_153_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_391 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_154_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_154_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_397 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_155_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_155_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_399 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_156_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_156_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_157_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_157_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_403 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_158_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_158_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_405 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_159_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_159_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_407 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_160_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_160_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_161_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_161_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_415 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_162_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_162_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_163_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_163_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_419 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_164_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_164_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_421 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_165_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_165_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_423 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_166_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_166_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_167_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_167_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_427 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_168_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_168_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_169_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_169_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_435 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_170_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_170_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_437 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_171_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_171_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_439 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_172_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_172_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_173_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_173_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_443 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_174_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_174_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_445 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_175_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_175_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_451 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_176_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_176_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_453 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_177_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_177_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_455 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_178_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_178_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_179_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_179_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_459 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_180_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_180_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_461 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_181_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_181_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_463 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_182_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_182_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_469 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_183_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_183_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_471 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_184_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_184_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_185_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_185_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_475 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_186_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_186_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_477 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_187_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_187_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_479 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_188_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_188_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_189_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_189_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_487 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_190_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_190_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_191_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_191_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_491 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_192_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_192_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_493 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_193_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_193_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_495 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_194_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_194_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_195_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_195_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_499 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_196_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_196_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_197_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_197_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_507 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_198_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_198_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_509 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_199_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_199_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_511 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_200_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_200_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_201_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_201_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_515 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_202_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_202_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_517 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_203_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_203_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_523 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_204_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_204_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_525 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_205_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_205_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_527 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_206_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_206_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_207_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_207_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_531 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_208_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_208_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_533 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_209_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_209_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_535 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_210_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_210_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_541 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_211_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_211_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_543 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_212_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_212_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_213_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_213_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_547 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_214_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_214_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_549 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_215_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_215_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_551 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_216_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_216_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_217_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_217_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_559 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_218_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_218_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_219_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_219_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_563 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_220_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_220_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_565 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_221_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_221_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_567 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_222_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_222_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_223_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_223_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_224_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_224_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_224_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_225_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_225_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[22], chanx_left_in[71]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size3 mux_bottom_track_35 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[24], chanx_left_in[75]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_bottom_out[17]));

	mux_tree_tapbuf_size3 mux_bottom_track_51 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[34], chanx_left_in[107]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_bottom_out[25]));

	mux_tree_tapbuf_size3 mux_bottom_track_53 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[36], chanx_left_in[111]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_bottom_out[26]));

	mux_tree_tapbuf_size3 mux_bottom_track_69 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[46], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_bottom_out[34]));

	mux_tree_tapbuf_size3 mux_bottom_track_71 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[48], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_bottom_out[35]));

	mux_tree_tapbuf_size3 mux_bottom_track_87 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[58], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_bottom_out[43]));

	mux_tree_tapbuf_size3 mux_bottom_track_89 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[60], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size3 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[70], chanx_left_in[215]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size3 mux_bottom_track_107 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[72], chanx_left_in[219]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_bottom_out[53]));

	mux_tree_tapbuf_size3 mux_bottom_track_123 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[82], chanx_left_in[251]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_bottom_out[61]));

	mux_tree_tapbuf_size3 mux_bottom_track_125 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[84], chanx_left_in[255]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_bottom_out[62]));

	mux_tree_tapbuf_size3 mux_bottom_track_141 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[94], chanx_left_in[284]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_bottom_out[70]));

	mux_tree_tapbuf_size3 mux_bottom_track_143 (
		.in({chanx_right_in[282], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_bottom_out[71]));

	mux_tree_tapbuf_size3 mux_bottom_track_159 (
		.in({chanx_right_in[272], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[106]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_bottom_out[79]));

	mux_tree_tapbuf_size3 mux_bottom_track_161 (
		.in({chanx_right_in[270], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[108]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size3 mux_bottom_track_177 (
		.in({chanx_right_in[260], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[118]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size3 mux_bottom_track_179 (
		.in({chanx_right_in[258], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[120]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_bottom_out[89]));

	mux_tree_tapbuf_size3 mux_bottom_track_195 (
		.in({chanx_right_in[248], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_bottom_out[97]));

	mux_tree_tapbuf_size3 mux_bottom_track_197 (
		.in({chanx_right_in[246], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_bottom_out[98]));

	mux_tree_tapbuf_size3 mux_bottom_track_213 (
		.in({chanx_right_in[236], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_bottom_out[106]));

	mux_tree_tapbuf_size3 mux_bottom_track_215 (
		.in({chanx_right_in[234], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_bottom_out[107]));

	mux_tree_tapbuf_size3 mux_bottom_track_231 (
		.in({chanx_right_in[224], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_bottom_out[115]));

	mux_tree_tapbuf_size3 mux_bottom_track_233 (
		.in({chanx_right_in[222], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size3 mux_bottom_track_249 (
		.in({chanx_right_in[212], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size3 mux_bottom_track_251 (
		.in({chanx_right_in[210], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_bottom_out[125]));

	mux_tree_tapbuf_size3 mux_bottom_track_267 (
		.in({chanx_right_in[200], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_bottom_out[133]));

	mux_tree_tapbuf_size3 mux_bottom_track_269 (
		.in({chanx_right_in[198], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_bottom_out[134]));

	mux_tree_tapbuf_size3 mux_bottom_track_285 (
		.in({chanx_right_in[188], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[190]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_bottom_out[142]));

	mux_tree_tapbuf_size3 mux_bottom_track_287 (
		.in({chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_bottom_out[143]));

	mux_tree_tapbuf_size3 mux_bottom_track_303 (
		.in({chanx_right_in[176], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[202]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_bottom_out[151]));

	mux_tree_tapbuf_size3 mux_bottom_track_305 (
		.in({chanx_right_in[174], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[204]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size3 mux_bottom_track_321 (
		.in({chanx_right_in[164], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[214]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size3 mux_bottom_track_323 (
		.in({chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[216]}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_bottom_out[161]));

	mux_tree_tapbuf_size3 mux_bottom_track_339 (
		.in({chanx_right_in[152], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[226]}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_bottom_out[169]));

	mux_tree_tapbuf_size3 mux_bottom_track_341 (
		.in({chanx_right_in[150], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[228]}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_bottom_out[170]));

	mux_tree_tapbuf_size3 mux_bottom_track_357 (
		.in({chanx_right_in[140], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[238]}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_bottom_out[178]));

	mux_tree_tapbuf_size3 mux_bottom_track_359 (
		.in({chanx_right_in[138], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[240]}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_bottom_out[179]));

	mux_tree_tapbuf_size3 mux_bottom_track_375 (
		.in({chanx_right_in[128], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[250]}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chany_bottom_out[187]));

	mux_tree_tapbuf_size3 mux_bottom_track_377 (
		.in({chanx_right_in[126], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[252]}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size3 mux_bottom_track_393 (
		.in({chanx_right_in[116], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[262]}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chany_bottom_out[196]));

	mux_tree_tapbuf_size3 mux_bottom_track_395 (
		.in({chanx_right_in[114], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[264]}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chany_bottom_out[197]));

	mux_tree_tapbuf_size3 mux_bottom_track_411 (
		.in({chanx_right_in[104], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[274]}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chany_bottom_out[205]));

	mux_tree_tapbuf_size3 mux_bottom_track_413 (
		.in({chanx_right_in[102], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[276]}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chany_bottom_out[206]));

	mux_tree_tapbuf_size3 mux_bottom_track_429 (
		.in({chanx_right_in[92], chanx_right_in[279], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chany_bottom_out[214]));

	mux_tree_tapbuf_size3 mux_bottom_track_431 (
		.in({chanx_right_in[90], chanx_right_in[275], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chany_bottom_out[215]));

	mux_tree_tapbuf_size3 mux_bottom_track_447 (
		.in({chanx_right_in[80], chanx_right_in[243], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chany_bottom_out[223]));

	mux_tree_tapbuf_size3 mux_bottom_track_449 (
		.in({chanx_right_in[78], chanx_right_in[239], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chany_bottom_out[224]));

	mux_tree_tapbuf_size3 mux_bottom_track_465 (
		.in({chanx_right_in[68], chanx_right_in[207], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chany_bottom_out[232]));

	mux_tree_tapbuf_size3 mux_bottom_track_467 (
		.in({chanx_right_in[66], chanx_right_in[203], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chany_bottom_out[233]));

	mux_tree_tapbuf_size3 mux_bottom_track_483 (
		.in({chanx_right_in[56], chanx_right_in[171], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chany_bottom_out[241]));

	mux_tree_tapbuf_size3 mux_bottom_track_485 (
		.in({chanx_right_in[54], chanx_right_in[167], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chany_bottom_out[242]));

	mux_tree_tapbuf_size3 mux_bottom_track_501 (
		.in({chanx_right_in[44], chanx_right_in[135], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chany_bottom_out[250]));

	mux_tree_tapbuf_size3 mux_bottom_track_503 (
		.in({chanx_right_in[42], chanx_right_in[131], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chany_bottom_out[251]));

	mux_tree_tapbuf_size3 mux_bottom_track_519 (
		.in({chanx_right_in[32], chanx_right_in[99], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chany_bottom_out[259]));

	mux_tree_tapbuf_size3 mux_bottom_track_521 (
		.in({chanx_right_in[30], chanx_right_in[95], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chany_bottom_out[260]));

	mux_tree_tapbuf_size3 mux_bottom_track_537 (
		.in({chanx_right_in[20], chanx_right_in[63], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chany_bottom_out[268]));

	mux_tree_tapbuf_size3 mux_bottom_track_539 (
		.in({chanx_right_in[18], chanx_right_in[59], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chany_bottom_out[269]));

	mux_tree_tapbuf_size3 mux_bottom_track_555 (
		.in({chanx_right_in[8], chanx_right_in[27], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chany_bottom_out[277]));

	mux_tree_tapbuf_size3 mux_bottom_track_557 (
		.in({chanx_right_in[6], chanx_right_in[23], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chany_bottom_out[278]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_213 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_215 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_231 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_251 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_267 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_269 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_285 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_287 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_303 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_323 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_339 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_341 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_357 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_359 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_375 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_395 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_411 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_413 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_429 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_431 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_447 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_467 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_483 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_485 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_501 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_503 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_519 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_539 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_555 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_bottom_track_557 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_1__18_ -----

//----- Default net type -----
`default_nettype wire



