//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: router]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 13:25:01 2024
//-------------------------------------------
// ----- BEGIN Grid Verilog module: grid_router -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for grid_router -----
module grid_router(reset,
                   clk,
                   top_width_0_height_0_subtile_0__pin_reset_0_,
                   top_width_0_height_0_subtile_0__pin_router_address_3_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_1_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_5_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_9_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_13_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_17_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_21_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_25_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_29_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_33_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_37_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_41_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_45_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_49_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_53_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_57_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_61_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_65_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_69_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_73_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_77_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_81_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_85_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_89_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_93_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_97_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_101_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_105_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_109_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_113_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_117_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_121_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_125_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_129_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_133_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_137_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_141_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_145_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_149_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_153_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_157_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_161_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_165_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_169_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_173_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_177_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_181_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_185_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_189_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_193_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_197_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_201_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_205_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_209_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_213_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_217_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_221_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_225_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_229_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_233_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_237_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_241_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_245_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_249_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_253_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_257_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_261_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_265_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_269_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_273_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_277_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_281_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_285_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_289_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_293_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_297_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_301_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_305_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_309_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_313_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_317_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_321_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_325_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_329_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_333_,
                   top_width_0_height_0_subtile_0__pin_channel_in_ip_337_,
                   top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_,
                   top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_,
                   top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_,
                   top_width_0_height_0_subtile_0__pin_clk_0_,
                   right_width_0_height_0_subtile_0__pin_router_address_0_,
                   right_width_0_height_0_subtile_0__pin_router_address_4_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_2_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_6_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_10_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_14_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_18_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_22_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_26_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_30_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_34_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_38_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_42_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_46_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_50_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_54_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_58_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_62_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_66_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_70_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_74_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_78_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_82_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_86_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_90_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_94_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_98_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_102_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_106_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_110_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_114_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_118_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_122_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_126_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_130_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_134_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_138_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_142_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_146_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_150_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_154_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_158_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_162_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_166_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_170_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_174_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_178_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_182_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_186_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_190_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_194_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_198_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_202_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_206_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_210_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_214_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_218_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_222_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_226_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_230_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_234_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_238_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_242_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_246_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_250_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_254_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_258_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_262_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_266_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_270_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_274_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_278_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_282_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_286_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_290_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_294_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_298_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_302_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_306_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_310_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_314_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_318_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_322_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_326_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_330_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_334_,
                   right_width_0_height_0_subtile_0__pin_channel_in_ip_338_,
                   right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_,
                   right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_,
                   bottom_width_0_height_0_subtile_0__pin_router_address_1_,
                   bottom_width_0_height_0_subtile_0__pin_router_address_5_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_,
                   bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_,
                   bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_,
                   bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_,
                   left_width_0_height_0_subtile_0__pin_router_address_2_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_0_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_4_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_8_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_12_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_16_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_20_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_24_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_28_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_32_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_36_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_40_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_44_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_48_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_52_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_56_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_60_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_64_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_68_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_72_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_76_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_80_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_84_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_88_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_92_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_96_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_100_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_104_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_108_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_112_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_116_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_120_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_124_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_128_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_132_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_136_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_140_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_144_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_148_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_152_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_156_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_160_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_164_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_168_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_172_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_176_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_180_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_184_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_188_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_192_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_196_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_200_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_204_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_208_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_212_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_216_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_220_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_224_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_228_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_232_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_236_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_240_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_244_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_248_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_252_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_256_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_260_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_264_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_268_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_272_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_276_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_280_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_284_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_288_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_292_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_296_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_300_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_304_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_308_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_312_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_316_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_320_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_324_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_328_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_332_,
                   left_width_0_height_0_subtile_0__pin_channel_in_ip_336_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_2_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_6_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_10_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_14_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_18_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_22_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_26_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_30_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_34_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_38_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_42_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_46_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_50_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_54_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_58_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_62_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_66_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_70_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_74_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_78_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_82_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_86_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_90_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_94_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_98_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_102_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_106_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_110_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_114_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_118_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_122_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_126_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_130_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_134_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_138_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_142_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_146_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_150_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_154_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_158_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_162_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_166_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_170_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_174_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_178_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_182_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_186_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_190_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_194_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_198_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_202_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_206_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_210_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_214_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_218_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_222_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_226_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_230_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_234_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_238_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_242_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_246_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_250_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_254_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_258_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_262_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_266_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_270_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_274_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_278_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_282_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_286_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_290_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_294_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_298_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_302_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_306_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_310_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_314_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_318_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_322_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_326_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_330_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_334_,
                   top_width_0_height_0_subtile_0__pin_channel_out_op_338_,
                   top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_,
                   top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_,
                   right_width_0_height_0_subtile_0__pin_error_0_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_3_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_7_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_11_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_15_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_19_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_23_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_27_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_31_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_35_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_39_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_43_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_47_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_51_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_55_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_59_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_63_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_67_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_71_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_75_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_79_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_83_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_87_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_91_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_95_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_99_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_103_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_107_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_111_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_115_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_119_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_123_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_127_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_131_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_135_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_139_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_143_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_147_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_151_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_155_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_159_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_163_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_167_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_171_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_175_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_179_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_183_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_187_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_191_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_195_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_199_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_203_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_207_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_211_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_215_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_219_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_223_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_227_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_231_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_235_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_239_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_243_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_247_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_251_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_255_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_259_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_263_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_267_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_271_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_275_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_279_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_283_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_287_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_291_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_295_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_299_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_303_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_307_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_311_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_315_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_319_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_323_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_327_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_331_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_335_,
                   right_width_0_height_0_subtile_0__pin_channel_out_op_339_,
                   right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_,
                   right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_,
                   bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_,
                   bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_,
                   bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_,
                   bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_1_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_5_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_9_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_13_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_17_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_21_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_25_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_29_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_33_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_37_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_41_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_45_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_49_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_53_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_57_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_61_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_65_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_69_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_73_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_77_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_81_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_85_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_89_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_93_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_97_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_101_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_105_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_109_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_113_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_117_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_121_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_125_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_129_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_133_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_137_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_141_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_145_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_149_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_153_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_157_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_161_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_165_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_169_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_173_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_177_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_181_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_185_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_189_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_193_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_197_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_201_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_205_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_209_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_213_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_217_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_221_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_225_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_229_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_233_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_237_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_241_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_245_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_249_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_253_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_257_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_261_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_265_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_269_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_273_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_277_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_281_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_285_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_289_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_293_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_297_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_301_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_305_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_309_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_313_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_317_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_321_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_325_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_329_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_333_,
                   left_width_0_height_0_subtile_0__pin_channel_out_op_337_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_,
                   left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_);
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_reset_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_router_address_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_33_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_37_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_41_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_45_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_49_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_53_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_57_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_61_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_65_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_69_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_73_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_77_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_81_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_85_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_89_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_93_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_97_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_101_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_105_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_109_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_113_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_117_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_121_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_125_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_129_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_133_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_137_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_141_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_145_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_149_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_153_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_157_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_161_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_165_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_169_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_173_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_177_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_181_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_185_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_189_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_193_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_197_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_201_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_205_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_209_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_213_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_217_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_221_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_225_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_229_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_233_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_237_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_241_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_245_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_249_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_253_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_257_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_261_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_265_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_269_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_273_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_277_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_281_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_285_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_289_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_293_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_297_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_301_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_305_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_309_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_313_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_317_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_321_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_325_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_329_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_333_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_channel_in_ip_337_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_router_address_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_router_address_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_router_address_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_router_address_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_router_address_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_20_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_24_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_28_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_32_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_36_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_40_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_44_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_48_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_52_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_56_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_60_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_64_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_68_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_72_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_76_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_80_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_84_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_88_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_92_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_96_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_100_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_104_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_108_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_112_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_116_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_120_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_124_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_128_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_132_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_136_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_140_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_144_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_148_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_152_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_156_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_160_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_164_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_168_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_172_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_176_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_180_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_184_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_188_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_192_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_196_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_200_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_204_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_208_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_212_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_216_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_220_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_224_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_228_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_232_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_236_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_240_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_244_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_248_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_252_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_256_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_260_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_264_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_268_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_272_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_276_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_280_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_284_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_288_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_292_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_296_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_300_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_304_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_308_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_312_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_316_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_320_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_324_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_328_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_332_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_channel_in_ip_336_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_error_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_router_mode_router_ logical_tile_router_mode_router__0 (
		.reset(reset),
		.clk(clk),
		.router_reset(top_width_0_height_0_subtile_0__pin_reset_0_),
		.router_router_address({right_width_0_height_0_subtile_0__pin_router_address_0_, bottom_width_0_height_0_subtile_0__pin_router_address_1_, left_width_0_height_0_subtile_0__pin_router_address_2_, top_width_0_height_0_subtile_0__pin_router_address_3_, right_width_0_height_0_subtile_0__pin_router_address_4_, bottom_width_0_height_0_subtile_0__pin_router_address_5_}),
		.router_channel_in_ip({left_width_0_height_0_subtile_0__pin_channel_in_ip_0_, top_width_0_height_0_subtile_0__pin_channel_in_ip_1_, right_width_0_height_0_subtile_0__pin_channel_in_ip_2_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_, left_width_0_height_0_subtile_0__pin_channel_in_ip_4_, top_width_0_height_0_subtile_0__pin_channel_in_ip_5_, right_width_0_height_0_subtile_0__pin_channel_in_ip_6_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_, left_width_0_height_0_subtile_0__pin_channel_in_ip_8_, top_width_0_height_0_subtile_0__pin_channel_in_ip_9_, right_width_0_height_0_subtile_0__pin_channel_in_ip_10_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_, left_width_0_height_0_subtile_0__pin_channel_in_ip_12_, top_width_0_height_0_subtile_0__pin_channel_in_ip_13_, right_width_0_height_0_subtile_0__pin_channel_in_ip_14_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_, left_width_0_height_0_subtile_0__pin_channel_in_ip_16_, top_width_0_height_0_subtile_0__pin_channel_in_ip_17_, right_width_0_height_0_subtile_0__pin_channel_in_ip_18_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_, left_width_0_height_0_subtile_0__pin_channel_in_ip_20_, top_width_0_height_0_subtile_0__pin_channel_in_ip_21_, right_width_0_height_0_subtile_0__pin_channel_in_ip_22_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_, left_width_0_height_0_subtile_0__pin_channel_in_ip_24_, top_width_0_height_0_subtile_0__pin_channel_in_ip_25_, right_width_0_height_0_subtile_0__pin_channel_in_ip_26_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_, left_width_0_height_0_subtile_0__pin_channel_in_ip_28_, top_width_0_height_0_subtile_0__pin_channel_in_ip_29_, right_width_0_height_0_subtile_0__pin_channel_in_ip_30_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_, left_width_0_height_0_subtile_0__pin_channel_in_ip_32_, top_width_0_height_0_subtile_0__pin_channel_in_ip_33_, right_width_0_height_0_subtile_0__pin_channel_in_ip_34_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_, left_width_0_height_0_subtile_0__pin_channel_in_ip_36_, top_width_0_height_0_subtile_0__pin_channel_in_ip_37_, right_width_0_height_0_subtile_0__pin_channel_in_ip_38_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_, left_width_0_height_0_subtile_0__pin_channel_in_ip_40_, top_width_0_height_0_subtile_0__pin_channel_in_ip_41_, right_width_0_height_0_subtile_0__pin_channel_in_ip_42_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_, left_width_0_height_0_subtile_0__pin_channel_in_ip_44_, top_width_0_height_0_subtile_0__pin_channel_in_ip_45_, right_width_0_height_0_subtile_0__pin_channel_in_ip_46_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_, left_width_0_height_0_subtile_0__pin_channel_in_ip_48_, top_width_0_height_0_subtile_0__pin_channel_in_ip_49_, right_width_0_height_0_subtile_0__pin_channel_in_ip_50_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_, left_width_0_height_0_subtile_0__pin_channel_in_ip_52_, top_width_0_height_0_subtile_0__pin_channel_in_ip_53_, right_width_0_height_0_subtile_0__pin_channel_in_ip_54_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_, left_width_0_height_0_subtile_0__pin_channel_in_ip_56_, top_width_0_height_0_subtile_0__pin_channel_in_ip_57_, right_width_0_height_0_subtile_0__pin_channel_in_ip_58_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_, left_width_0_height_0_subtile_0__pin_channel_in_ip_60_, top_width_0_height_0_subtile_0__pin_channel_in_ip_61_, right_width_0_height_0_subtile_0__pin_channel_in_ip_62_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_, left_width_0_height_0_subtile_0__pin_channel_in_ip_64_, top_width_0_height_0_subtile_0__pin_channel_in_ip_65_, right_width_0_height_0_subtile_0__pin_channel_in_ip_66_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_, left_width_0_height_0_subtile_0__pin_channel_in_ip_68_, top_width_0_height_0_subtile_0__pin_channel_in_ip_69_, right_width_0_height_0_subtile_0__pin_channel_in_ip_70_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_, left_width_0_height_0_subtile_0__pin_channel_in_ip_72_, top_width_0_height_0_subtile_0__pin_channel_in_ip_73_, right_width_0_height_0_subtile_0__pin_channel_in_ip_74_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_, left_width_0_height_0_subtile_0__pin_channel_in_ip_76_, top_width_0_height_0_subtile_0__pin_channel_in_ip_77_, right_width_0_height_0_subtile_0__pin_channel_in_ip_78_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_, left_width_0_height_0_subtile_0__pin_channel_in_ip_80_, top_width_0_height_0_subtile_0__pin_channel_in_ip_81_, right_width_0_height_0_subtile_0__pin_channel_in_ip_82_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_, left_width_0_height_0_subtile_0__pin_channel_in_ip_84_, top_width_0_height_0_subtile_0__pin_channel_in_ip_85_, right_width_0_height_0_subtile_0__pin_channel_in_ip_86_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_, left_width_0_height_0_subtile_0__pin_channel_in_ip_88_, top_width_0_height_0_subtile_0__pin_channel_in_ip_89_, right_width_0_height_0_subtile_0__pin_channel_in_ip_90_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_, left_width_0_height_0_subtile_0__pin_channel_in_ip_92_, top_width_0_height_0_subtile_0__pin_channel_in_ip_93_, right_width_0_height_0_subtile_0__pin_channel_in_ip_94_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_, left_width_0_height_0_subtile_0__pin_channel_in_ip_96_, top_width_0_height_0_subtile_0__pin_channel_in_ip_97_, right_width_0_height_0_subtile_0__pin_channel_in_ip_98_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_, left_width_0_height_0_subtile_0__pin_channel_in_ip_100_, top_width_0_height_0_subtile_0__pin_channel_in_ip_101_, right_width_0_height_0_subtile_0__pin_channel_in_ip_102_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_, left_width_0_height_0_subtile_0__pin_channel_in_ip_104_, top_width_0_height_0_subtile_0__pin_channel_in_ip_105_, right_width_0_height_0_subtile_0__pin_channel_in_ip_106_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_, left_width_0_height_0_subtile_0__pin_channel_in_ip_108_, top_width_0_height_0_subtile_0__pin_channel_in_ip_109_, right_width_0_height_0_subtile_0__pin_channel_in_ip_110_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_, left_width_0_height_0_subtile_0__pin_channel_in_ip_112_, top_width_0_height_0_subtile_0__pin_channel_in_ip_113_, right_width_0_height_0_subtile_0__pin_channel_in_ip_114_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_, left_width_0_height_0_subtile_0__pin_channel_in_ip_116_, top_width_0_height_0_subtile_0__pin_channel_in_ip_117_, right_width_0_height_0_subtile_0__pin_channel_in_ip_118_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_, left_width_0_height_0_subtile_0__pin_channel_in_ip_120_, top_width_0_height_0_subtile_0__pin_channel_in_ip_121_, right_width_0_height_0_subtile_0__pin_channel_in_ip_122_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_, left_width_0_height_0_subtile_0__pin_channel_in_ip_124_, top_width_0_height_0_subtile_0__pin_channel_in_ip_125_, right_width_0_height_0_subtile_0__pin_channel_in_ip_126_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_, left_width_0_height_0_subtile_0__pin_channel_in_ip_128_, top_width_0_height_0_subtile_0__pin_channel_in_ip_129_, right_width_0_height_0_subtile_0__pin_channel_in_ip_130_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_, left_width_0_height_0_subtile_0__pin_channel_in_ip_132_, top_width_0_height_0_subtile_0__pin_channel_in_ip_133_, right_width_0_height_0_subtile_0__pin_channel_in_ip_134_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_, left_width_0_height_0_subtile_0__pin_channel_in_ip_136_, top_width_0_height_0_subtile_0__pin_channel_in_ip_137_, right_width_0_height_0_subtile_0__pin_channel_in_ip_138_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_, left_width_0_height_0_subtile_0__pin_channel_in_ip_140_, top_width_0_height_0_subtile_0__pin_channel_in_ip_141_, right_width_0_height_0_subtile_0__pin_channel_in_ip_142_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_, left_width_0_height_0_subtile_0__pin_channel_in_ip_144_, top_width_0_height_0_subtile_0__pin_channel_in_ip_145_, right_width_0_height_0_subtile_0__pin_channel_in_ip_146_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_, left_width_0_height_0_subtile_0__pin_channel_in_ip_148_, top_width_0_height_0_subtile_0__pin_channel_in_ip_149_, right_width_0_height_0_subtile_0__pin_channel_in_ip_150_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_, left_width_0_height_0_subtile_0__pin_channel_in_ip_152_, top_width_0_height_0_subtile_0__pin_channel_in_ip_153_, right_width_0_height_0_subtile_0__pin_channel_in_ip_154_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_, left_width_0_height_0_subtile_0__pin_channel_in_ip_156_, top_width_0_height_0_subtile_0__pin_channel_in_ip_157_, right_width_0_height_0_subtile_0__pin_channel_in_ip_158_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_, left_width_0_height_0_subtile_0__pin_channel_in_ip_160_, top_width_0_height_0_subtile_0__pin_channel_in_ip_161_, right_width_0_height_0_subtile_0__pin_channel_in_ip_162_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_, left_width_0_height_0_subtile_0__pin_channel_in_ip_164_, top_width_0_height_0_subtile_0__pin_channel_in_ip_165_, right_width_0_height_0_subtile_0__pin_channel_in_ip_166_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_, left_width_0_height_0_subtile_0__pin_channel_in_ip_168_, top_width_0_height_0_subtile_0__pin_channel_in_ip_169_, right_width_0_height_0_subtile_0__pin_channel_in_ip_170_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_, left_width_0_height_0_subtile_0__pin_channel_in_ip_172_, top_width_0_height_0_subtile_0__pin_channel_in_ip_173_, right_width_0_height_0_subtile_0__pin_channel_in_ip_174_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_, left_width_0_height_0_subtile_0__pin_channel_in_ip_176_, top_width_0_height_0_subtile_0__pin_channel_in_ip_177_, right_width_0_height_0_subtile_0__pin_channel_in_ip_178_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_, left_width_0_height_0_subtile_0__pin_channel_in_ip_180_, top_width_0_height_0_subtile_0__pin_channel_in_ip_181_, right_width_0_height_0_subtile_0__pin_channel_in_ip_182_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_, left_width_0_height_0_subtile_0__pin_channel_in_ip_184_, top_width_0_height_0_subtile_0__pin_channel_in_ip_185_, right_width_0_height_0_subtile_0__pin_channel_in_ip_186_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_, left_width_0_height_0_subtile_0__pin_channel_in_ip_188_, top_width_0_height_0_subtile_0__pin_channel_in_ip_189_, right_width_0_height_0_subtile_0__pin_channel_in_ip_190_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_, left_width_0_height_0_subtile_0__pin_channel_in_ip_192_, top_width_0_height_0_subtile_0__pin_channel_in_ip_193_, right_width_0_height_0_subtile_0__pin_channel_in_ip_194_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_, left_width_0_height_0_subtile_0__pin_channel_in_ip_196_, top_width_0_height_0_subtile_0__pin_channel_in_ip_197_, right_width_0_height_0_subtile_0__pin_channel_in_ip_198_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_, left_width_0_height_0_subtile_0__pin_channel_in_ip_200_, top_width_0_height_0_subtile_0__pin_channel_in_ip_201_, right_width_0_height_0_subtile_0__pin_channel_in_ip_202_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_, left_width_0_height_0_subtile_0__pin_channel_in_ip_204_, top_width_0_height_0_subtile_0__pin_channel_in_ip_205_, right_width_0_height_0_subtile_0__pin_channel_in_ip_206_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_, left_width_0_height_0_subtile_0__pin_channel_in_ip_208_, top_width_0_height_0_subtile_0__pin_channel_in_ip_209_, right_width_0_height_0_subtile_0__pin_channel_in_ip_210_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_, left_width_0_height_0_subtile_0__pin_channel_in_ip_212_, top_width_0_height_0_subtile_0__pin_channel_in_ip_213_, right_width_0_height_0_subtile_0__pin_channel_in_ip_214_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_, left_width_0_height_0_subtile_0__pin_channel_in_ip_216_, top_width_0_height_0_subtile_0__pin_channel_in_ip_217_, right_width_0_height_0_subtile_0__pin_channel_in_ip_218_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_, left_width_0_height_0_subtile_0__pin_channel_in_ip_220_, top_width_0_height_0_subtile_0__pin_channel_in_ip_221_, right_width_0_height_0_subtile_0__pin_channel_in_ip_222_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_, left_width_0_height_0_subtile_0__pin_channel_in_ip_224_, top_width_0_height_0_subtile_0__pin_channel_in_ip_225_, right_width_0_height_0_subtile_0__pin_channel_in_ip_226_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_, left_width_0_height_0_subtile_0__pin_channel_in_ip_228_, top_width_0_height_0_subtile_0__pin_channel_in_ip_229_, right_width_0_height_0_subtile_0__pin_channel_in_ip_230_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_, left_width_0_height_0_subtile_0__pin_channel_in_ip_232_, top_width_0_height_0_subtile_0__pin_channel_in_ip_233_, right_width_0_height_0_subtile_0__pin_channel_in_ip_234_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_, left_width_0_height_0_subtile_0__pin_channel_in_ip_236_, top_width_0_height_0_subtile_0__pin_channel_in_ip_237_, right_width_0_height_0_subtile_0__pin_channel_in_ip_238_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_, left_width_0_height_0_subtile_0__pin_channel_in_ip_240_, top_width_0_height_0_subtile_0__pin_channel_in_ip_241_, right_width_0_height_0_subtile_0__pin_channel_in_ip_242_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_, left_width_0_height_0_subtile_0__pin_channel_in_ip_244_, top_width_0_height_0_subtile_0__pin_channel_in_ip_245_, right_width_0_height_0_subtile_0__pin_channel_in_ip_246_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_, left_width_0_height_0_subtile_0__pin_channel_in_ip_248_, top_width_0_height_0_subtile_0__pin_channel_in_ip_249_, right_width_0_height_0_subtile_0__pin_channel_in_ip_250_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_, left_width_0_height_0_subtile_0__pin_channel_in_ip_252_, top_width_0_height_0_subtile_0__pin_channel_in_ip_253_, right_width_0_height_0_subtile_0__pin_channel_in_ip_254_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_, left_width_0_height_0_subtile_0__pin_channel_in_ip_256_, top_width_0_height_0_subtile_0__pin_channel_in_ip_257_, right_width_0_height_0_subtile_0__pin_channel_in_ip_258_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_, left_width_0_height_0_subtile_0__pin_channel_in_ip_260_, top_width_0_height_0_subtile_0__pin_channel_in_ip_261_, right_width_0_height_0_subtile_0__pin_channel_in_ip_262_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_, left_width_0_height_0_subtile_0__pin_channel_in_ip_264_, top_width_0_height_0_subtile_0__pin_channel_in_ip_265_, right_width_0_height_0_subtile_0__pin_channel_in_ip_266_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_, left_width_0_height_0_subtile_0__pin_channel_in_ip_268_, top_width_0_height_0_subtile_0__pin_channel_in_ip_269_, right_width_0_height_0_subtile_0__pin_channel_in_ip_270_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_, left_width_0_height_0_subtile_0__pin_channel_in_ip_272_, top_width_0_height_0_subtile_0__pin_channel_in_ip_273_, right_width_0_height_0_subtile_0__pin_channel_in_ip_274_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_, left_width_0_height_0_subtile_0__pin_channel_in_ip_276_, top_width_0_height_0_subtile_0__pin_channel_in_ip_277_, right_width_0_height_0_subtile_0__pin_channel_in_ip_278_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_, left_width_0_height_0_subtile_0__pin_channel_in_ip_280_, top_width_0_height_0_subtile_0__pin_channel_in_ip_281_, right_width_0_height_0_subtile_0__pin_channel_in_ip_282_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_, left_width_0_height_0_subtile_0__pin_channel_in_ip_284_, top_width_0_height_0_subtile_0__pin_channel_in_ip_285_, right_width_0_height_0_subtile_0__pin_channel_in_ip_286_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_, left_width_0_height_0_subtile_0__pin_channel_in_ip_288_, top_width_0_height_0_subtile_0__pin_channel_in_ip_289_, right_width_0_height_0_subtile_0__pin_channel_in_ip_290_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_, left_width_0_height_0_subtile_0__pin_channel_in_ip_292_, top_width_0_height_0_subtile_0__pin_channel_in_ip_293_, right_width_0_height_0_subtile_0__pin_channel_in_ip_294_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_, left_width_0_height_0_subtile_0__pin_channel_in_ip_296_, top_width_0_height_0_subtile_0__pin_channel_in_ip_297_, right_width_0_height_0_subtile_0__pin_channel_in_ip_298_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_, left_width_0_height_0_subtile_0__pin_channel_in_ip_300_, top_width_0_height_0_subtile_0__pin_channel_in_ip_301_, right_width_0_height_0_subtile_0__pin_channel_in_ip_302_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_, left_width_0_height_0_subtile_0__pin_channel_in_ip_304_, top_width_0_height_0_subtile_0__pin_channel_in_ip_305_, right_width_0_height_0_subtile_0__pin_channel_in_ip_306_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_, left_width_0_height_0_subtile_0__pin_channel_in_ip_308_, top_width_0_height_0_subtile_0__pin_channel_in_ip_309_, right_width_0_height_0_subtile_0__pin_channel_in_ip_310_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_, left_width_0_height_0_subtile_0__pin_channel_in_ip_312_, top_width_0_height_0_subtile_0__pin_channel_in_ip_313_, right_width_0_height_0_subtile_0__pin_channel_in_ip_314_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_, left_width_0_height_0_subtile_0__pin_channel_in_ip_316_, top_width_0_height_0_subtile_0__pin_channel_in_ip_317_, right_width_0_height_0_subtile_0__pin_channel_in_ip_318_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_, left_width_0_height_0_subtile_0__pin_channel_in_ip_320_, top_width_0_height_0_subtile_0__pin_channel_in_ip_321_, right_width_0_height_0_subtile_0__pin_channel_in_ip_322_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_, left_width_0_height_0_subtile_0__pin_channel_in_ip_324_, top_width_0_height_0_subtile_0__pin_channel_in_ip_325_, right_width_0_height_0_subtile_0__pin_channel_in_ip_326_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_, left_width_0_height_0_subtile_0__pin_channel_in_ip_328_, top_width_0_height_0_subtile_0__pin_channel_in_ip_329_, right_width_0_height_0_subtile_0__pin_channel_in_ip_330_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_, left_width_0_height_0_subtile_0__pin_channel_in_ip_332_, top_width_0_height_0_subtile_0__pin_channel_in_ip_333_, right_width_0_height_0_subtile_0__pin_channel_in_ip_334_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_, left_width_0_height_0_subtile_0__pin_channel_in_ip_336_, top_width_0_height_0_subtile_0__pin_channel_in_ip_337_, right_width_0_height_0_subtile_0__pin_channel_in_ip_338_, bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_}),
		.router_flow_ctrl_in_op({left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_, top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_, right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_, bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_, left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_, top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_, right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_, bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_, left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_, top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_}),
		.router_clk(top_width_0_height_0_subtile_0__pin_clk_0_),
		.router_error(right_width_0_height_0_subtile_0__pin_error_0_),
		.router_channel_out_op({bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_width_0_height_0_subtile_0__pin_channel_out_op_302_, right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, left_width_0_height_0_subtile_0__pin_channel_out_op_305_, top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_width_0_height_0_subtile_0__pin_channel_out_op_310_, right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_width_0_height_0_subtile_0__pin_channel_out_op_314_, right_width_0_height_0_subtile_0__pin_channel_out_op_315_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, left_width_0_height_0_subtile_0__pin_channel_out_op_317_, top_width_0_height_0_subtile_0__pin_channel_out_op_318_, right_width_0_height_0_subtile_0__pin_channel_out_op_319_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, left_width_0_height_0_subtile_0__pin_channel_out_op_321_, top_width_0_height_0_subtile_0__pin_channel_out_op_322_, right_width_0_height_0_subtile_0__pin_channel_out_op_323_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, left_width_0_height_0_subtile_0__pin_channel_out_op_325_, top_width_0_height_0_subtile_0__pin_channel_out_op_326_, right_width_0_height_0_subtile_0__pin_channel_out_op_327_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, left_width_0_height_0_subtile_0__pin_channel_out_op_329_, top_width_0_height_0_subtile_0__pin_channel_out_op_330_, right_width_0_height_0_subtile_0__pin_channel_out_op_331_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, left_width_0_height_0_subtile_0__pin_channel_out_op_333_, top_width_0_height_0_subtile_0__pin_channel_out_op_334_, right_width_0_height_0_subtile_0__pin_channel_out_op_335_, bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, left_width_0_height_0_subtile_0__pin_channel_out_op_337_, top_width_0_height_0_subtile_0__pin_channel_out_op_338_, right_width_0_height_0_subtile_0__pin_channel_out_op_339_}),
		.router_flow_ctrl_out_ip({bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_}));

endmodule
// ----- END Verilog module for grid_router -----

//----- Default net type -----
`default_nettype wire



// ----- END Grid Verilog module: grid_router -----

