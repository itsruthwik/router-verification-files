//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Jul 24 20:28:26 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:479] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:104] cbx_1__0__0_chanx_left_out;
wire [0:104] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__10_ccff_tail;
wire [0:104] cbx_1__0__10_chanx_left_out;
wire [0:104] cbx_1__0__10_chanx_right_out;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__11_ccff_tail;
wire [0:104] cbx_1__0__11_chanx_left_out;
wire [0:104] cbx_1__0__11_chanx_right_out;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__12_ccff_tail;
wire [0:104] cbx_1__0__12_chanx_left_out;
wire [0:104] cbx_1__0__12_chanx_right_out;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__13_ccff_tail;
wire [0:104] cbx_1__0__13_chanx_left_out;
wire [0:104] cbx_1__0__13_chanx_right_out;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__14_ccff_tail;
wire [0:104] cbx_1__0__14_chanx_left_out;
wire [0:104] cbx_1__0__14_chanx_right_out;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__15_ccff_tail;
wire [0:104] cbx_1__0__15_chanx_left_out;
wire [0:104] cbx_1__0__15_chanx_right_out;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__16_ccff_tail;
wire [0:104] cbx_1__0__16_chanx_left_out;
wire [0:104] cbx_1__0__16_chanx_right_out;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__17_ccff_tail;
wire [0:104] cbx_1__0__17_chanx_left_out;
wire [0:104] cbx_1__0__17_chanx_right_out;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__18_ccff_tail;
wire [0:104] cbx_1__0__18_chanx_left_out;
wire [0:104] cbx_1__0__18_chanx_right_out;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__19_ccff_tail;
wire [0:104] cbx_1__0__19_chanx_left_out;
wire [0:104] cbx_1__0__19_chanx_right_out;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:104] cbx_1__0__1_chanx_left_out;
wire [0:104] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:104] cbx_1__0__2_chanx_left_out;
wire [0:104] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:104] cbx_1__0__3_chanx_left_out;
wire [0:104] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__4_ccff_tail;
wire [0:104] cbx_1__0__4_chanx_left_out;
wire [0:104] cbx_1__0__4_chanx_right_out;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__5_ccff_tail;
wire [0:104] cbx_1__0__5_chanx_left_out;
wire [0:104] cbx_1__0__5_chanx_right_out;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__6_ccff_tail;
wire [0:104] cbx_1__0__6_chanx_left_out;
wire [0:104] cbx_1__0__6_chanx_right_out;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__7_ccff_tail;
wire [0:104] cbx_1__0__7_chanx_left_out;
wire [0:104] cbx_1__0__7_chanx_right_out;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__8_ccff_tail;
wire [0:104] cbx_1__0__8_chanx_left_out;
wire [0:104] cbx_1__0__8_chanx_right_out;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__9_ccff_tail;
wire [0:104] cbx_1__0__9_chanx_left_out;
wire [0:104] cbx_1__0__9_chanx_right_out;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__0_ccff_tail;
wire [0:104] cbx_1__10__0_chanx_left_out;
wire [0:104] cbx_1__10__0_chanx_right_out;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__1_ccff_tail;
wire [0:104] cbx_1__10__1_chanx_left_out;
wire [0:104] cbx_1__10__1_chanx_right_out;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__2_ccff_tail;
wire [0:104] cbx_1__10__2_chanx_left_out;
wire [0:104] cbx_1__10__2_chanx_right_out;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__3_ccff_tail;
wire [0:104] cbx_1__10__3_chanx_left_out;
wire [0:104] cbx_1__10__3_chanx_right_out;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__4_ccff_tail;
wire [0:104] cbx_1__10__4_chanx_left_out;
wire [0:104] cbx_1__10__4_chanx_right_out;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__5_ccff_tail;
wire [0:104] cbx_1__10__5_chanx_left_out;
wire [0:104] cbx_1__10__5_chanx_right_out;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__6_ccff_tail;
wire [0:104] cbx_1__10__6_chanx_left_out;
wire [0:104] cbx_1__10__6_chanx_right_out;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__7_ccff_tail;
wire [0:104] cbx_1__10__7_chanx_left_out;
wire [0:104] cbx_1__10__7_chanx_right_out;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__8_ccff_tail;
wire [0:104] cbx_1__10__8_chanx_left_out;
wire [0:104] cbx_1__10__8_chanx_right_out;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__10__9_ccff_tail;
wire [0:104] cbx_1__10__9_chanx_left_out;
wire [0:104] cbx_1__10__9_chanx_right_out;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:104] cbx_1__2__0_chanx_left_out;
wire [0:104] cbx_1__2__0_chanx_right_out;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:104] cbx_1__2__1_chanx_left_out;
wire [0:104] cbx_1__2__1_chanx_right_out;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__2_ccff_tail;
wire [0:104] cbx_1__2__2_chanx_left_out;
wire [0:104] cbx_1__2__2_chanx_right_out;
wire [0:0] cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__3_ccff_tail;
wire [0:104] cbx_1__2__3_chanx_left_out;
wire [0:104] cbx_1__2__3_chanx_right_out;
wire [0:0] cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__4_ccff_tail;
wire [0:104] cbx_1__2__4_chanx_left_out;
wire [0:104] cbx_1__2__4_chanx_right_out;
wire [0:0] cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__5_ccff_tail;
wire [0:104] cbx_1__2__5_chanx_left_out;
wire [0:104] cbx_1__2__5_chanx_right_out;
wire [0:0] cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__6_ccff_tail;
wire [0:104] cbx_1__2__6_chanx_left_out;
wire [0:104] cbx_1__2__6_chanx_right_out;
wire [0:0] cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__7_ccff_tail;
wire [0:104] cbx_1__2__7_chanx_left_out;
wire [0:104] cbx_1__2__7_chanx_right_out;
wire [0:0] cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__8_ccff_tail;
wire [0:104] cbx_1__2__8_chanx_left_out;
wire [0:104] cbx_1__2__8_chanx_right_out;
wire [0:0] cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__2__9_ccff_tail;
wire [0:104] cbx_1__2__9_chanx_left_out;
wire [0:104] cbx_1__2__9_chanx_right_out;
wire [0:0] cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__0_ccff_tail;
wire [0:104] cbx_1__3__0_chanx_left_out;
wire [0:104] cbx_1__3__0_chanx_right_out;
wire [0:0] cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__10_ccff_tail;
wire [0:104] cbx_1__3__10_chanx_left_out;
wire [0:104] cbx_1__3__10_chanx_right_out;
wire [0:0] cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__11_ccff_tail;
wire [0:104] cbx_1__3__11_chanx_left_out;
wire [0:104] cbx_1__3__11_chanx_right_out;
wire [0:0] cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__12_ccff_tail;
wire [0:104] cbx_1__3__12_chanx_left_out;
wire [0:104] cbx_1__3__12_chanx_right_out;
wire [0:0] cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__13_ccff_tail;
wire [0:104] cbx_1__3__13_chanx_left_out;
wire [0:104] cbx_1__3__13_chanx_right_out;
wire [0:0] cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__14_ccff_tail;
wire [0:104] cbx_1__3__14_chanx_left_out;
wire [0:104] cbx_1__3__14_chanx_right_out;
wire [0:0] cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__15_ccff_tail;
wire [0:104] cbx_1__3__15_chanx_left_out;
wire [0:104] cbx_1__3__15_chanx_right_out;
wire [0:0] cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__16_ccff_tail;
wire [0:104] cbx_1__3__16_chanx_left_out;
wire [0:104] cbx_1__3__16_chanx_right_out;
wire [0:0] cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__17_ccff_tail;
wire [0:104] cbx_1__3__17_chanx_left_out;
wire [0:104] cbx_1__3__17_chanx_right_out;
wire [0:0] cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__18_ccff_tail;
wire [0:104] cbx_1__3__18_chanx_left_out;
wire [0:104] cbx_1__3__18_chanx_right_out;
wire [0:0] cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__19_ccff_tail;
wire [0:104] cbx_1__3__19_chanx_left_out;
wire [0:104] cbx_1__3__19_chanx_right_out;
wire [0:0] cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__1_ccff_tail;
wire [0:104] cbx_1__3__1_chanx_left_out;
wire [0:104] cbx_1__3__1_chanx_right_out;
wire [0:0] cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__20_ccff_tail;
wire [0:104] cbx_1__3__20_chanx_left_out;
wire [0:104] cbx_1__3__20_chanx_right_out;
wire [0:0] cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__21_ccff_tail;
wire [0:104] cbx_1__3__21_chanx_left_out;
wire [0:104] cbx_1__3__21_chanx_right_out;
wire [0:0] cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__22_ccff_tail;
wire [0:104] cbx_1__3__22_chanx_left_out;
wire [0:104] cbx_1__3__22_chanx_right_out;
wire [0:0] cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__23_ccff_tail;
wire [0:104] cbx_1__3__23_chanx_left_out;
wire [0:104] cbx_1__3__23_chanx_right_out;
wire [0:0] cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__24_ccff_tail;
wire [0:104] cbx_1__3__24_chanx_left_out;
wire [0:104] cbx_1__3__24_chanx_right_out;
wire [0:0] cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__25_ccff_tail;
wire [0:104] cbx_1__3__25_chanx_left_out;
wire [0:104] cbx_1__3__25_chanx_right_out;
wire [0:0] cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__26_ccff_tail;
wire [0:104] cbx_1__3__26_chanx_left_out;
wire [0:104] cbx_1__3__26_chanx_right_out;
wire [0:0] cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__27_ccff_tail;
wire [0:104] cbx_1__3__27_chanx_left_out;
wire [0:104] cbx_1__3__27_chanx_right_out;
wire [0:0] cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__28_ccff_tail;
wire [0:104] cbx_1__3__28_chanx_left_out;
wire [0:104] cbx_1__3__28_chanx_right_out;
wire [0:0] cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__29_ccff_tail;
wire [0:104] cbx_1__3__29_chanx_left_out;
wire [0:104] cbx_1__3__29_chanx_right_out;
wire [0:0] cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__2_ccff_tail;
wire [0:104] cbx_1__3__2_chanx_left_out;
wire [0:104] cbx_1__3__2_chanx_right_out;
wire [0:0] cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__30_ccff_tail;
wire [0:104] cbx_1__3__30_chanx_left_out;
wire [0:104] cbx_1__3__30_chanx_right_out;
wire [0:0] cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__31_ccff_tail;
wire [0:104] cbx_1__3__31_chanx_left_out;
wire [0:104] cbx_1__3__31_chanx_right_out;
wire [0:0] cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__32_ccff_tail;
wire [0:104] cbx_1__3__32_chanx_left_out;
wire [0:104] cbx_1__3__32_chanx_right_out;
wire [0:0] cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__33_ccff_tail;
wire [0:104] cbx_1__3__33_chanx_left_out;
wire [0:104] cbx_1__3__33_chanx_right_out;
wire [0:0] cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__34_ccff_tail;
wire [0:104] cbx_1__3__34_chanx_left_out;
wire [0:104] cbx_1__3__34_chanx_right_out;
wire [0:0] cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__35_ccff_tail;
wire [0:104] cbx_1__3__35_chanx_left_out;
wire [0:104] cbx_1__3__35_chanx_right_out;
wire [0:0] cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__36_ccff_tail;
wire [0:104] cbx_1__3__36_chanx_left_out;
wire [0:104] cbx_1__3__36_chanx_right_out;
wire [0:0] cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__37_ccff_tail;
wire [0:104] cbx_1__3__37_chanx_left_out;
wire [0:104] cbx_1__3__37_chanx_right_out;
wire [0:0] cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__38_ccff_tail;
wire [0:104] cbx_1__3__38_chanx_left_out;
wire [0:104] cbx_1__3__38_chanx_right_out;
wire [0:0] cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__39_ccff_tail;
wire [0:104] cbx_1__3__39_chanx_left_out;
wire [0:104] cbx_1__3__39_chanx_right_out;
wire [0:0] cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__3_ccff_tail;
wire [0:104] cbx_1__3__3_chanx_left_out;
wire [0:104] cbx_1__3__3_chanx_right_out;
wire [0:0] cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__40_ccff_tail;
wire [0:104] cbx_1__3__40_chanx_left_out;
wire [0:104] cbx_1__3__40_chanx_right_out;
wire [0:0] cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__41_ccff_tail;
wire [0:104] cbx_1__3__41_chanx_left_out;
wire [0:104] cbx_1__3__41_chanx_right_out;
wire [0:0] cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__42_ccff_tail;
wire [0:104] cbx_1__3__42_chanx_left_out;
wire [0:104] cbx_1__3__42_chanx_right_out;
wire [0:0] cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__43_ccff_tail;
wire [0:104] cbx_1__3__43_chanx_left_out;
wire [0:104] cbx_1__3__43_chanx_right_out;
wire [0:0] cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__44_ccff_tail;
wire [0:104] cbx_1__3__44_chanx_left_out;
wire [0:104] cbx_1__3__44_chanx_right_out;
wire [0:0] cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__45_ccff_tail;
wire [0:104] cbx_1__3__45_chanx_left_out;
wire [0:104] cbx_1__3__45_chanx_right_out;
wire [0:0] cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__46_ccff_tail;
wire [0:104] cbx_1__3__46_chanx_left_out;
wire [0:104] cbx_1__3__46_chanx_right_out;
wire [0:0] cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__47_ccff_tail;
wire [0:104] cbx_1__3__47_chanx_left_out;
wire [0:104] cbx_1__3__47_chanx_right_out;
wire [0:0] cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__48_ccff_tail;
wire [0:104] cbx_1__3__48_chanx_left_out;
wire [0:104] cbx_1__3__48_chanx_right_out;
wire [0:0] cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__49_ccff_tail;
wire [0:104] cbx_1__3__49_chanx_left_out;
wire [0:104] cbx_1__3__49_chanx_right_out;
wire [0:0] cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__4_ccff_tail;
wire [0:104] cbx_1__3__4_chanx_left_out;
wire [0:104] cbx_1__3__4_chanx_right_out;
wire [0:0] cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__50_ccff_tail;
wire [0:104] cbx_1__3__50_chanx_left_out;
wire [0:104] cbx_1__3__50_chanx_right_out;
wire [0:0] cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__51_ccff_tail;
wire [0:104] cbx_1__3__51_chanx_left_out;
wire [0:104] cbx_1__3__51_chanx_right_out;
wire [0:0] cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__52_ccff_tail;
wire [0:104] cbx_1__3__52_chanx_left_out;
wire [0:104] cbx_1__3__52_chanx_right_out;
wire [0:0] cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__53_ccff_tail;
wire [0:104] cbx_1__3__53_chanx_left_out;
wire [0:104] cbx_1__3__53_chanx_right_out;
wire [0:0] cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__54_ccff_tail;
wire [0:104] cbx_1__3__54_chanx_left_out;
wire [0:104] cbx_1__3__54_chanx_right_out;
wire [0:0] cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__55_ccff_tail;
wire [0:104] cbx_1__3__55_chanx_left_out;
wire [0:104] cbx_1__3__55_chanx_right_out;
wire [0:0] cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__56_ccff_tail;
wire [0:104] cbx_1__3__56_chanx_left_out;
wire [0:104] cbx_1__3__56_chanx_right_out;
wire [0:0] cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__57_ccff_tail;
wire [0:104] cbx_1__3__57_chanx_left_out;
wire [0:104] cbx_1__3__57_chanx_right_out;
wire [0:0] cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__58_ccff_tail;
wire [0:104] cbx_1__3__58_chanx_left_out;
wire [0:104] cbx_1__3__58_chanx_right_out;
wire [0:0] cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__59_ccff_tail;
wire [0:104] cbx_1__3__59_chanx_left_out;
wire [0:104] cbx_1__3__59_chanx_right_out;
wire [0:0] cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__5_ccff_tail;
wire [0:104] cbx_1__3__5_chanx_left_out;
wire [0:104] cbx_1__3__5_chanx_right_out;
wire [0:0] cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__60_ccff_tail;
wire [0:104] cbx_1__3__60_chanx_left_out;
wire [0:104] cbx_1__3__60_chanx_right_out;
wire [0:0] cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__61_ccff_tail;
wire [0:104] cbx_1__3__61_chanx_left_out;
wire [0:104] cbx_1__3__61_chanx_right_out;
wire [0:0] cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__62_ccff_tail;
wire [0:104] cbx_1__3__62_chanx_left_out;
wire [0:104] cbx_1__3__62_chanx_right_out;
wire [0:0] cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__63_ccff_tail;
wire [0:104] cbx_1__3__63_chanx_left_out;
wire [0:104] cbx_1__3__63_chanx_right_out;
wire [0:0] cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__64_ccff_tail;
wire [0:104] cbx_1__3__64_chanx_left_out;
wire [0:104] cbx_1__3__64_chanx_right_out;
wire [0:0] cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__65_ccff_tail;
wire [0:104] cbx_1__3__65_chanx_left_out;
wire [0:104] cbx_1__3__65_chanx_right_out;
wire [0:0] cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__6_ccff_tail;
wire [0:104] cbx_1__3__6_chanx_left_out;
wire [0:104] cbx_1__3__6_chanx_right_out;
wire [0:0] cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__7_ccff_tail;
wire [0:104] cbx_1__3__7_chanx_left_out;
wire [0:104] cbx_1__3__7_chanx_right_out;
wire [0:0] cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__8_ccff_tail;
wire [0:104] cbx_1__3__8_chanx_left_out;
wire [0:104] cbx_1__3__8_chanx_right_out;
wire [0:0] cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__9_ccff_tail;
wire [0:104] cbx_1__3__9_chanx_left_out;
wire [0:104] cbx_1__3__9_chanx_right_out;
wire [0:0] cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_6__5__0_ccff_tail;
wire [0:104] cbx_6__5__0_chanx_left_out;
wire [0:104] cbx_6__5__0_chanx_right_out;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_6__5__1_ccff_tail;
wire [0:104] cbx_6__5__1_chanx_left_out;
wire [0:104] cbx_6__5__1_chanx_right_out;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
wire [0:0] cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_6__6__0_ccff_tail;
wire [0:104] cbx_6__6__0_chanx_left_out;
wire [0:104] cbx_6__6__0_chanx_right_out;
wire [0:0] cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_;
wire [0:0] cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_;
wire [0:0] cbx_6__6__1_ccff_tail;
wire [0:104] cbx_6__6__1_chanx_left_out;
wire [0:104] cbx_6__6__1_chanx_right_out;
wire [0:0] cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:104] cby_0__1__0_chany_bottom_out;
wire [0:104] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__10_ccff_tail;
wire [0:104] cby_0__1__10_chany_bottom_out;
wire [0:104] cby_0__1__10_chany_top_out;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__11_ccff_tail;
wire [0:104] cby_0__1__11_chany_bottom_out;
wire [0:104] cby_0__1__11_chany_top_out;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__12_ccff_tail;
wire [0:104] cby_0__1__12_chany_bottom_out;
wire [0:104] cby_0__1__12_chany_top_out;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__13_ccff_tail;
wire [0:104] cby_0__1__13_chany_bottom_out;
wire [0:104] cby_0__1__13_chany_top_out;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__14_ccff_tail;
wire [0:104] cby_0__1__14_chany_bottom_out;
wire [0:104] cby_0__1__14_chany_top_out;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__15_ccff_tail;
wire [0:104] cby_0__1__15_chany_bottom_out;
wire [0:104] cby_0__1__15_chany_top_out;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__16_ccff_tail;
wire [0:104] cby_0__1__16_chany_bottom_out;
wire [0:104] cby_0__1__16_chany_top_out;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__17_ccff_tail;
wire [0:104] cby_0__1__17_chany_bottom_out;
wire [0:104] cby_0__1__17_chany_top_out;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__18_ccff_tail;
wire [0:104] cby_0__1__18_chany_bottom_out;
wire [0:104] cby_0__1__18_chany_top_out;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__19_ccff_tail;
wire [0:104] cby_0__1__19_chany_bottom_out;
wire [0:104] cby_0__1__19_chany_top_out;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:104] cby_0__1__1_chany_bottom_out;
wire [0:104] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__20_ccff_tail;
wire [0:104] cby_0__1__20_chany_bottom_out;
wire [0:104] cby_0__1__20_chany_top_out;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__21_ccff_tail;
wire [0:104] cby_0__1__21_chany_bottom_out;
wire [0:104] cby_0__1__21_chany_top_out;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__21_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__21_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:104] cby_0__1__2_chany_bottom_out;
wire [0:104] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:104] cby_0__1__3_chany_bottom_out;
wire [0:104] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__4_ccff_tail;
wire [0:104] cby_0__1__4_chany_bottom_out;
wire [0:104] cby_0__1__4_chany_top_out;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__5_ccff_tail;
wire [0:104] cby_0__1__5_chany_bottom_out;
wire [0:104] cby_0__1__5_chany_top_out;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__6_ccff_tail;
wire [0:104] cby_0__1__6_chany_bottom_out;
wire [0:104] cby_0__1__6_chany_top_out;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__7_ccff_tail;
wire [0:104] cby_0__1__7_chany_bottom_out;
wire [0:104] cby_0__1__7_chany_top_out;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__8_ccff_tail;
wire [0:104] cby_0__1__8_chany_bottom_out;
wire [0:104] cby_0__1__8_chany_top_out;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__9_ccff_tail;
wire [0:104] cby_0__1__9_chany_bottom_out;
wire [0:104] cby_0__1__9_chany_top_out;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__0_ccff_tail;
wire [0:104] cby_0__3__0_chany_bottom_out;
wire [0:104] cby_0__3__0_chany_top_out;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__1_ccff_tail;
wire [0:104] cby_0__3__1_chany_bottom_out;
wire [0:104] cby_0__3__1_chany_top_out;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__2_ccff_tail;
wire [0:104] cby_0__3__2_chany_bottom_out;
wire [0:104] cby_0__3__2_chany_top_out;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__3_ccff_tail;
wire [0:104] cby_0__3__3_chany_bottom_out;
wire [0:104] cby_0__3__3_chany_top_out;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__4_ccff_tail;
wire [0:104] cby_0__3__4_chany_bottom_out;
wire [0:104] cby_0__3__4_chany_top_out;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__5_ccff_tail;
wire [0:104] cby_0__3__5_chany_bottom_out;
wire [0:104] cby_0__3__5_chany_top_out;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__6_ccff_tail;
wire [0:104] cby_0__3__6_chany_bottom_out;
wire [0:104] cby_0__3__6_chany_top_out;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__3__7_ccff_tail;
wire [0:104] cby_0__3__7_chany_bottom_out;
wire [0:104] cby_0__3__7_chany_top_out;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__3__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_10__3__0_ccff_tail;
wire [0:104] cby_10__3__0_chany_bottom_out;
wire [0:104] cby_10__3__0_chany_top_out;
wire [0:0] cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__1_ccff_tail;
wire [0:104] cby_10__3__1_chany_bottom_out;
wire [0:104] cby_10__3__1_chany_top_out;
wire [0:0] cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__2_ccff_tail;
wire [0:104] cby_10__3__2_chany_bottom_out;
wire [0:104] cby_10__3__2_chany_top_out;
wire [0:0] cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__3_ccff_tail;
wire [0:104] cby_10__3__3_chany_bottom_out;
wire [0:104] cby_10__3__3_chany_top_out;
wire [0:0] cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__4_ccff_tail;
wire [0:104] cby_10__3__4_chany_bottom_out;
wire [0:104] cby_10__3__4_chany_top_out;
wire [0:0] cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__5_ccff_tail;
wire [0:104] cby_10__3__5_chany_bottom_out;
wire [0:104] cby_10__3__5_chany_top_out;
wire [0:0] cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__3__6_ccff_tail;
wire [0:104] cby_10__3__6_chany_bottom_out;
wire [0:104] cby_10__3__6_chany_top_out;
wire [0:0] cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__3__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_10__6__0_ccff_tail;
wire [0:104] cby_10__6__0_chany_bottom_out;
wire [0:104] cby_10__6__0_chany_top_out;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_10__6__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_1__3__0_ccff_tail;
wire [0:104] cby_1__3__0_chany_bottom_out;
wire [0:104] cby_1__3__0_chany_top_out;
wire [0:0] cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__10_ccff_tail;
wire [0:104] cby_1__3__10_chany_bottom_out;
wire [0:104] cby_1__3__10_chany_top_out;
wire [0:0] cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__11_ccff_tail;
wire [0:104] cby_1__3__11_chany_bottom_out;
wire [0:104] cby_1__3__11_chany_top_out;
wire [0:0] cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__12_ccff_tail;
wire [0:104] cby_1__3__12_chany_bottom_out;
wire [0:104] cby_1__3__12_chany_top_out;
wire [0:0] cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__13_ccff_tail;
wire [0:104] cby_1__3__13_chany_bottom_out;
wire [0:104] cby_1__3__13_chany_top_out;
wire [0:0] cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__14_ccff_tail;
wire [0:104] cby_1__3__14_chany_bottom_out;
wire [0:104] cby_1__3__14_chany_top_out;
wire [0:0] cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__15_ccff_tail;
wire [0:104] cby_1__3__15_chany_bottom_out;
wire [0:104] cby_1__3__15_chany_top_out;
wire [0:0] cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__16_ccff_tail;
wire [0:104] cby_1__3__16_chany_bottom_out;
wire [0:104] cby_1__3__16_chany_top_out;
wire [0:0] cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__17_ccff_tail;
wire [0:104] cby_1__3__17_chany_bottom_out;
wire [0:104] cby_1__3__17_chany_top_out;
wire [0:0] cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__18_ccff_tail;
wire [0:104] cby_1__3__18_chany_bottom_out;
wire [0:104] cby_1__3__18_chany_top_out;
wire [0:0] cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__19_ccff_tail;
wire [0:104] cby_1__3__19_chany_bottom_out;
wire [0:104] cby_1__3__19_chany_top_out;
wire [0:0] cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__1_ccff_tail;
wire [0:104] cby_1__3__1_chany_bottom_out;
wire [0:104] cby_1__3__1_chany_top_out;
wire [0:0] cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__20_ccff_tail;
wire [0:104] cby_1__3__20_chany_bottom_out;
wire [0:104] cby_1__3__20_chany_top_out;
wire [0:0] cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__21_ccff_tail;
wire [0:104] cby_1__3__21_chany_bottom_out;
wire [0:104] cby_1__3__21_chany_top_out;
wire [0:0] cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__22_ccff_tail;
wire [0:104] cby_1__3__22_chany_bottom_out;
wire [0:104] cby_1__3__22_chany_top_out;
wire [0:0] cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__23_ccff_tail;
wire [0:104] cby_1__3__23_chany_bottom_out;
wire [0:104] cby_1__3__23_chany_top_out;
wire [0:0] cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__24_ccff_tail;
wire [0:104] cby_1__3__24_chany_bottom_out;
wire [0:104] cby_1__3__24_chany_top_out;
wire [0:0] cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__25_ccff_tail;
wire [0:104] cby_1__3__25_chany_bottom_out;
wire [0:104] cby_1__3__25_chany_top_out;
wire [0:0] cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__26_ccff_tail;
wire [0:104] cby_1__3__26_chany_bottom_out;
wire [0:104] cby_1__3__26_chany_top_out;
wire [0:0] cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__27_ccff_tail;
wire [0:104] cby_1__3__27_chany_bottom_out;
wire [0:104] cby_1__3__27_chany_top_out;
wire [0:0] cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__28_ccff_tail;
wire [0:104] cby_1__3__28_chany_bottom_out;
wire [0:104] cby_1__3__28_chany_top_out;
wire [0:0] cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__29_ccff_tail;
wire [0:104] cby_1__3__29_chany_bottom_out;
wire [0:104] cby_1__3__29_chany_top_out;
wire [0:0] cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__2_ccff_tail;
wire [0:104] cby_1__3__2_chany_bottom_out;
wire [0:104] cby_1__3__2_chany_top_out;
wire [0:0] cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__30_ccff_tail;
wire [0:104] cby_1__3__30_chany_bottom_out;
wire [0:104] cby_1__3__30_chany_top_out;
wire [0:0] cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__31_ccff_tail;
wire [0:104] cby_1__3__31_chany_bottom_out;
wire [0:104] cby_1__3__31_chany_top_out;
wire [0:0] cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__32_ccff_tail;
wire [0:104] cby_1__3__32_chany_bottom_out;
wire [0:104] cby_1__3__32_chany_top_out;
wire [0:0] cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__33_ccff_tail;
wire [0:104] cby_1__3__33_chany_bottom_out;
wire [0:104] cby_1__3__33_chany_top_out;
wire [0:0] cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__34_ccff_tail;
wire [0:104] cby_1__3__34_chany_bottom_out;
wire [0:104] cby_1__3__34_chany_top_out;
wire [0:0] cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__35_ccff_tail;
wire [0:104] cby_1__3__35_chany_bottom_out;
wire [0:104] cby_1__3__35_chany_top_out;
wire [0:0] cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__36_ccff_tail;
wire [0:104] cby_1__3__36_chany_bottom_out;
wire [0:104] cby_1__3__36_chany_top_out;
wire [0:0] cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__37_ccff_tail;
wire [0:104] cby_1__3__37_chany_bottom_out;
wire [0:104] cby_1__3__37_chany_top_out;
wire [0:0] cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__38_ccff_tail;
wire [0:104] cby_1__3__38_chany_bottom_out;
wire [0:104] cby_1__3__38_chany_top_out;
wire [0:0] cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__39_ccff_tail;
wire [0:104] cby_1__3__39_chany_bottom_out;
wire [0:104] cby_1__3__39_chany_top_out;
wire [0:0] cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__3_ccff_tail;
wire [0:104] cby_1__3__3_chany_bottom_out;
wire [0:104] cby_1__3__3_chany_top_out;
wire [0:0] cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__40_ccff_tail;
wire [0:104] cby_1__3__40_chany_bottom_out;
wire [0:104] cby_1__3__40_chany_top_out;
wire [0:0] cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__41_ccff_tail;
wire [0:104] cby_1__3__41_chany_bottom_out;
wire [0:104] cby_1__3__41_chany_top_out;
wire [0:0] cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__42_ccff_tail;
wire [0:104] cby_1__3__42_chany_bottom_out;
wire [0:104] cby_1__3__42_chany_top_out;
wire [0:0] cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__43_ccff_tail;
wire [0:104] cby_1__3__43_chany_bottom_out;
wire [0:104] cby_1__3__43_chany_top_out;
wire [0:0] cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__44_ccff_tail;
wire [0:104] cby_1__3__44_chany_bottom_out;
wire [0:104] cby_1__3__44_chany_top_out;
wire [0:0] cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__45_ccff_tail;
wire [0:104] cby_1__3__45_chany_bottom_out;
wire [0:104] cby_1__3__45_chany_top_out;
wire [0:0] cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__46_ccff_tail;
wire [0:104] cby_1__3__46_chany_bottom_out;
wire [0:104] cby_1__3__46_chany_top_out;
wire [0:0] cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__47_ccff_tail;
wire [0:104] cby_1__3__47_chany_bottom_out;
wire [0:104] cby_1__3__47_chany_top_out;
wire [0:0] cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__48_ccff_tail;
wire [0:104] cby_1__3__48_chany_bottom_out;
wire [0:104] cby_1__3__48_chany_top_out;
wire [0:0] cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__49_ccff_tail;
wire [0:104] cby_1__3__49_chany_bottom_out;
wire [0:104] cby_1__3__49_chany_top_out;
wire [0:0] cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__4_ccff_tail;
wire [0:104] cby_1__3__4_chany_bottom_out;
wire [0:104] cby_1__3__4_chany_top_out;
wire [0:0] cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__50_ccff_tail;
wire [0:104] cby_1__3__50_chany_bottom_out;
wire [0:104] cby_1__3__50_chany_top_out;
wire [0:0] cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__51_ccff_tail;
wire [0:104] cby_1__3__51_chany_bottom_out;
wire [0:104] cby_1__3__51_chany_top_out;
wire [0:0] cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__52_ccff_tail;
wire [0:104] cby_1__3__52_chany_bottom_out;
wire [0:104] cby_1__3__52_chany_top_out;
wire [0:0] cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__53_ccff_tail;
wire [0:104] cby_1__3__53_chany_bottom_out;
wire [0:104] cby_1__3__53_chany_top_out;
wire [0:0] cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__54_ccff_tail;
wire [0:104] cby_1__3__54_chany_bottom_out;
wire [0:104] cby_1__3__54_chany_top_out;
wire [0:0] cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__55_ccff_tail;
wire [0:104] cby_1__3__55_chany_bottom_out;
wire [0:104] cby_1__3__55_chany_top_out;
wire [0:0] cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__56_ccff_tail;
wire [0:104] cby_1__3__56_chany_bottom_out;
wire [0:104] cby_1__3__56_chany_top_out;
wire [0:0] cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__57_ccff_tail;
wire [0:104] cby_1__3__57_chany_bottom_out;
wire [0:104] cby_1__3__57_chany_top_out;
wire [0:0] cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__58_ccff_tail;
wire [0:104] cby_1__3__58_chany_bottom_out;
wire [0:104] cby_1__3__58_chany_top_out;
wire [0:0] cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__59_ccff_tail;
wire [0:104] cby_1__3__59_chany_bottom_out;
wire [0:104] cby_1__3__59_chany_top_out;
wire [0:0] cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__5_ccff_tail;
wire [0:104] cby_1__3__5_chany_bottom_out;
wire [0:104] cby_1__3__5_chany_top_out;
wire [0:0] cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__60_ccff_tail;
wire [0:104] cby_1__3__60_chany_bottom_out;
wire [0:104] cby_1__3__60_chany_top_out;
wire [0:0] cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__61_ccff_tail;
wire [0:104] cby_1__3__61_chany_bottom_out;
wire [0:104] cby_1__3__61_chany_top_out;
wire [0:0] cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__62_ccff_tail;
wire [0:104] cby_1__3__62_chany_bottom_out;
wire [0:104] cby_1__3__62_chany_top_out;
wire [0:0] cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__63_ccff_tail;
wire [0:104] cby_1__3__63_chany_bottom_out;
wire [0:104] cby_1__3__63_chany_top_out;
wire [0:0] cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__64_ccff_tail;
wire [0:104] cby_1__3__64_chany_bottom_out;
wire [0:104] cby_1__3__64_chany_top_out;
wire [0:0] cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__65_ccff_tail;
wire [0:104] cby_1__3__65_chany_bottom_out;
wire [0:104] cby_1__3__65_chany_top_out;
wire [0:0] cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__66_ccff_tail;
wire [0:104] cby_1__3__66_chany_bottom_out;
wire [0:104] cby_1__3__66_chany_top_out;
wire [0:0] cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__67_ccff_tail;
wire [0:104] cby_1__3__67_chany_bottom_out;
wire [0:104] cby_1__3__67_chany_top_out;
wire [0:0] cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__68_ccff_tail;
wire [0:104] cby_1__3__68_chany_bottom_out;
wire [0:104] cby_1__3__68_chany_top_out;
wire [0:0] cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__6_ccff_tail;
wire [0:104] cby_1__3__6_chany_bottom_out;
wire [0:104] cby_1__3__6_chany_top_out;
wire [0:0] cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__7_ccff_tail;
wire [0:104] cby_1__3__7_chany_bottom_out;
wire [0:104] cby_1__3__7_chany_top_out;
wire [0:0] cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__8_ccff_tail;
wire [0:104] cby_1__3__8_chany_bottom_out;
wire [0:104] cby_1__3__8_chany_top_out;
wire [0:0] cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__3__9_ccff_tail;
wire [0:104] cby_1__3__9_chany_bottom_out;
wire [0:104] cby_1__3__9_chany_top_out;
wire [0:0] cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_5__6__0_ccff_tail;
wire [0:104] cby_5__6__0_chany_bottom_out;
wire [0:104] cby_5__6__0_chany_top_out;
wire [0:0] cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_5__6__1_ccff_tail;
wire [0:104] cby_5__6__1_chany_bottom_out;
wire [0:104] cby_5__6__1_chany_top_out;
wire [0:0] cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_;
wire [0:0] cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_;
wire [0:0] cby_6__6__0_ccff_tail;
wire [0:104] cby_6__6__0_chany_bottom_out;
wire [0:104] cby_6__6__0_chany_top_out;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_;
wire [0:0] cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_;
wire [0:0] cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_10__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_20_ccff_tail;
wire [0:0] grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_21_ccff_tail;
wire [0:0] grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_22_ccff_tail;
wire [0:0] grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_23_ccff_tail;
wire [0:0] grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_24_ccff_tail;
wire [0:0] grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_25_ccff_tail;
wire [0:0] grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_26_ccff_tail;
wire [0:0] grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_27_ccff_tail;
wire [0:0] grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_28_ccff_tail;
wire [0:0] grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_29_ccff_tail;
wire [0:0] grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_2__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_30_ccff_tail;
wire [0:0] grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_31_ccff_tail;
wire [0:0] grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_32_ccff_tail;
wire [0:0] grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_33_ccff_tail;
wire [0:0] grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_34_ccff_tail;
wire [0:0] grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_35_ccff_tail;
wire [0:0] grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_36_ccff_tail;
wire [0:0] grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_37_ccff_tail;
wire [0:0] grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_38_ccff_tail;
wire [0:0] grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_39_ccff_tail;
wire [0:0] grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3_ccff_tail;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_40_ccff_tail;
wire [0:0] grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_41_ccff_tail;
wire [0:0] grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_42_ccff_tail;
wire [0:0] grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_43_ccff_tail;
wire [0:0] grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_44_ccff_tail;
wire [0:0] grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_45_ccff_tail;
wire [0:0] grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_46_ccff_tail;
wire [0:0] grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_47_ccff_tail;
wire [0:0] grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_48_ccff_tail;
wire [0:0] grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_49_ccff_tail;
wire [0:0] grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_50_ccff_tail;
wire [0:0] grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_51_ccff_tail;
wire [0:0] grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_52_ccff_tail;
wire [0:0] grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_53_ccff_tail;
wire [0:0] grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_54_ccff_tail;
wire [0:0] grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_55_ccff_tail;
wire [0:0] grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_56_ccff_tail;
wire [0:0] grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_57_ccff_tail;
wire [0:0] grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_58_ccff_tail;
wire [0:0] grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_59_ccff_tail;
wire [0:0] grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_60_ccff_tail;
wire [0:0] grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_61_ccff_tail;
wire [0:0] grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_62_ccff_tail;
wire [0:0] grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_63_ccff_tail;
wire [0:0] grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_64_ccff_tail;
wire [0:0] grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_65_ccff_tail;
wire [0:0] grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_66_ccff_tail;
wire [0:0] grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_67_ccff_tail;
wire [0:0] grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_68_ccff_tail;
wire [0:0] grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_69_ccff_tail;
wire [0:0] grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_6__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_70_ccff_tail;
wire [0:0] grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_71_ccff_tail;
wire [0:0] grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_72_ccff_tail;
wire [0:0] grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_73_ccff_tail;
wire [0:0] grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_74_ccff_tail;
wire [0:0] grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_75_ccff_tail;
wire [0:0] grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_76_ccff_tail;
wire [0:0] grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_77_ccff_tail;
wire [0:0] grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_8__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_9__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_0_ccff_tail;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_10_ccff_tail;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_10_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_10_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_10_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_11_ccff_tail;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_11_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_11_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_11_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_12_ccff_tail;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_12_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_12_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_12_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_13_ccff_tail;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_13_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_13_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_13_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_14_ccff_tail;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_14_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_14_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_14_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_15_ccff_tail;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_15_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_15_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_15_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_16_ccff_tail;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_16_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_16_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_16_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_17_ccff_tail;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_17_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_17_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_17_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_18_ccff_tail;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_18_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_18_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_18_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_19_ccff_tail;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_19_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_19_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_19_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_1_ccff_tail;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_2_ccff_tail;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_2_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_2_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_3_ccff_tail;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_3_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_3_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_4_ccff_tail;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_4_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_4_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_4_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_5_ccff_tail;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_5_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_5_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_5_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_6_ccff_tail;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_6_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_6_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_6_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_7_ccff_tail;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_7_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_7_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_7_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_8_ccff_tail;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_8_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_8_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_8_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_9_ccff_tail;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_9_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_9_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_9_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_ccff_tail;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_ccff_tail;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_ccff_tail;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_ccff_tail;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_ccff_tail;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_ccff_tail;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_2_ccff_tail;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_3_ccff_tail;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_4_ccff_tail;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_5_ccff_tail;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_6_ccff_tail;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_7_ccff_tail;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_8_ccff_tail;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_9_ccff_tail;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_2_ccff_tail;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_3_ccff_tail;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_4_ccff_tail;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_5_ccff_tail;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_6_ccff_tail;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_7_ccff_tail;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_8_ccff_tail;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_9_ccff_tail;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_2_ccff_tail;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_3_ccff_tail;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_4_ccff_tail;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_5_ccff_tail;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_6_ccff_tail;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_7_ccff_tail;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_8_ccff_tail;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_9_ccff_tail;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_10__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_;
wire [0:0] grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:104] sb_0__0__0_chanx_right_out;
wire [0:104] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__10__0_ccff_tail;
wire [0:104] sb_0__10__0_chanx_right_out;
wire [0:104] sb_0__10__0_chany_bottom_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:104] sb_0__1__0_chanx_right_out;
wire [0:104] sb_0__1__0_chany_bottom_out;
wire [0:104] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:104] sb_0__2__0_chanx_right_out;
wire [0:104] sb_0__2__0_chany_bottom_out;
wire [0:104] sb_0__2__0_chany_top_out;
wire [0:0] sb_0__3__0_ccff_tail;
wire [0:104] sb_0__3__0_chanx_right_out;
wire [0:104] sb_0__3__0_chany_bottom_out;
wire [0:104] sb_0__3__0_chany_top_out;
wire [0:0] sb_0__3__1_ccff_tail;
wire [0:104] sb_0__3__1_chanx_right_out;
wire [0:104] sb_0__3__1_chany_bottom_out;
wire [0:104] sb_0__3__1_chany_top_out;
wire [0:0] sb_0__3__2_ccff_tail;
wire [0:104] sb_0__3__2_chanx_right_out;
wire [0:104] sb_0__3__2_chany_bottom_out;
wire [0:104] sb_0__3__2_chany_top_out;
wire [0:0] sb_0__3__3_ccff_tail;
wire [0:104] sb_0__3__3_chanx_right_out;
wire [0:104] sb_0__3__3_chany_bottom_out;
wire [0:104] sb_0__3__3_chany_top_out;
wire [0:0] sb_0__3__4_ccff_tail;
wire [0:104] sb_0__3__4_chanx_right_out;
wire [0:104] sb_0__3__4_chany_bottom_out;
wire [0:104] sb_0__3__4_chany_top_out;
wire [0:0] sb_0__3__5_ccff_tail;
wire [0:104] sb_0__3__5_chanx_right_out;
wire [0:104] sb_0__3__5_chany_bottom_out;
wire [0:104] sb_0__3__5_chany_top_out;
wire [0:0] sb_0__3__6_ccff_tail;
wire [0:104] sb_0__3__6_chanx_right_out;
wire [0:104] sb_0__3__6_chany_bottom_out;
wire [0:104] sb_0__3__6_chany_top_out;
wire [0:0] sb_10__0__0_ccff_tail;
wire [0:104] sb_10__0__0_chanx_left_out;
wire [0:104] sb_10__0__0_chany_top_out;
wire [0:0] sb_10__10__0_ccff_tail;
wire [0:104] sb_10__10__0_chanx_left_out;
wire [0:104] sb_10__10__0_chany_bottom_out;
wire [0:0] sb_10__1__0_ccff_tail;
wire [0:104] sb_10__1__0_chanx_left_out;
wire [0:104] sb_10__1__0_chany_bottom_out;
wire [0:104] sb_10__1__0_chany_top_out;
wire [0:0] sb_10__2__0_ccff_tail;
wire [0:104] sb_10__2__0_chanx_left_out;
wire [0:104] sb_10__2__0_chany_bottom_out;
wire [0:104] sb_10__2__0_chany_top_out;
wire [0:0] sb_10__3__0_ccff_tail;
wire [0:104] sb_10__3__0_chanx_left_out;
wire [0:104] sb_10__3__0_chany_bottom_out;
wire [0:104] sb_10__3__0_chany_top_out;
wire [0:0] sb_10__3__1_ccff_tail;
wire [0:104] sb_10__3__1_chanx_left_out;
wire [0:104] sb_10__3__1_chany_bottom_out;
wire [0:104] sb_10__3__1_chany_top_out;
wire [0:0] sb_10__3__2_ccff_tail;
wire [0:104] sb_10__3__2_chanx_left_out;
wire [0:104] sb_10__3__2_chany_bottom_out;
wire [0:104] sb_10__3__2_chany_top_out;
wire [0:0] sb_10__3__3_ccff_tail;
wire [0:104] sb_10__3__3_chanx_left_out;
wire [0:104] sb_10__3__3_chany_bottom_out;
wire [0:104] sb_10__3__3_chany_top_out;
wire [0:0] sb_10__3__4_ccff_tail;
wire [0:104] sb_10__3__4_chanx_left_out;
wire [0:104] sb_10__3__4_chany_bottom_out;
wire [0:104] sb_10__3__4_chany_top_out;
wire [0:0] sb_10__5__0_ccff_tail;
wire [0:104] sb_10__5__0_chanx_left_out;
wire [0:104] sb_10__5__0_chany_bottom_out;
wire [0:104] sb_10__5__0_chany_top_out;
wire [0:0] sb_10__6__0_ccff_tail;
wire [0:104] sb_10__6__0_chanx_left_out;
wire [0:104] sb_10__6__0_chany_bottom_out;
wire [0:104] sb_10__6__0_chany_top_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:104] sb_1__0__0_chanx_left_out;
wire [0:104] sb_1__0__0_chanx_right_out;
wire [0:104] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:104] sb_1__0__1_chanx_left_out;
wire [0:104] sb_1__0__1_chanx_right_out;
wire [0:104] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:104] sb_1__0__2_chanx_left_out;
wire [0:104] sb_1__0__2_chanx_right_out;
wire [0:104] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__0__3_ccff_tail;
wire [0:104] sb_1__0__3_chanx_left_out;
wire [0:104] sb_1__0__3_chanx_right_out;
wire [0:104] sb_1__0__3_chany_top_out;
wire [0:0] sb_1__0__4_ccff_tail;
wire [0:104] sb_1__0__4_chanx_left_out;
wire [0:104] sb_1__0__4_chanx_right_out;
wire [0:104] sb_1__0__4_chany_top_out;
wire [0:0] sb_1__0__5_ccff_tail;
wire [0:104] sb_1__0__5_chanx_left_out;
wire [0:104] sb_1__0__5_chanx_right_out;
wire [0:104] sb_1__0__5_chany_top_out;
wire [0:0] sb_1__0__6_ccff_tail;
wire [0:104] sb_1__0__6_chanx_left_out;
wire [0:104] sb_1__0__6_chanx_right_out;
wire [0:104] sb_1__0__6_chany_top_out;
wire [0:0] sb_1__0__7_ccff_tail;
wire [0:104] sb_1__0__7_chanx_left_out;
wire [0:104] sb_1__0__7_chanx_right_out;
wire [0:104] sb_1__0__7_chany_top_out;
wire [0:0] sb_1__0__8_ccff_tail;
wire [0:104] sb_1__0__8_chanx_left_out;
wire [0:104] sb_1__0__8_chanx_right_out;
wire [0:104] sb_1__0__8_chany_top_out;
wire [0:0] sb_1__10__0_ccff_tail;
wire [0:104] sb_1__10__0_chanx_left_out;
wire [0:104] sb_1__10__0_chanx_right_out;
wire [0:104] sb_1__10__0_chany_bottom_out;
wire [0:0] sb_1__10__1_ccff_tail;
wire [0:104] sb_1__10__1_chanx_left_out;
wire [0:104] sb_1__10__1_chanx_right_out;
wire [0:104] sb_1__10__1_chany_bottom_out;
wire [0:0] sb_1__10__2_ccff_tail;
wire [0:104] sb_1__10__2_chanx_left_out;
wire [0:104] sb_1__10__2_chanx_right_out;
wire [0:104] sb_1__10__2_chany_bottom_out;
wire [0:0] sb_1__10__3_ccff_tail;
wire [0:104] sb_1__10__3_chanx_left_out;
wire [0:104] sb_1__10__3_chanx_right_out;
wire [0:104] sb_1__10__3_chany_bottom_out;
wire [0:0] sb_1__10__4_ccff_tail;
wire [0:104] sb_1__10__4_chanx_left_out;
wire [0:104] sb_1__10__4_chanx_right_out;
wire [0:104] sb_1__10__4_chany_bottom_out;
wire [0:0] sb_1__10__5_ccff_tail;
wire [0:104] sb_1__10__5_chanx_left_out;
wire [0:104] sb_1__10__5_chanx_right_out;
wire [0:104] sb_1__10__5_chany_bottom_out;
wire [0:0] sb_1__10__6_ccff_tail;
wire [0:104] sb_1__10__6_chanx_left_out;
wire [0:104] sb_1__10__6_chanx_right_out;
wire [0:104] sb_1__10__6_chany_bottom_out;
wire [0:0] sb_1__10__7_ccff_tail;
wire [0:104] sb_1__10__7_chanx_left_out;
wire [0:104] sb_1__10__7_chanx_right_out;
wire [0:104] sb_1__10__7_chany_bottom_out;
wire [0:0] sb_1__10__8_ccff_tail;
wire [0:104] sb_1__10__8_chanx_left_out;
wire [0:104] sb_1__10__8_chanx_right_out;
wire [0:104] sb_1__10__8_chany_bottom_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:104] sb_1__1__0_chanx_left_out;
wire [0:104] sb_1__1__0_chanx_right_out;
wire [0:104] sb_1__1__0_chany_bottom_out;
wire [0:104] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:104] sb_1__1__1_chanx_left_out;
wire [0:104] sb_1__1__1_chanx_right_out;
wire [0:104] sb_1__1__1_chany_bottom_out;
wire [0:104] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__1__2_ccff_tail;
wire [0:104] sb_1__1__2_chanx_left_out;
wire [0:104] sb_1__1__2_chanx_right_out;
wire [0:104] sb_1__1__2_chany_bottom_out;
wire [0:104] sb_1__1__2_chany_top_out;
wire [0:0] sb_1__1__3_ccff_tail;
wire [0:104] sb_1__1__3_chanx_left_out;
wire [0:104] sb_1__1__3_chanx_right_out;
wire [0:104] sb_1__1__3_chany_bottom_out;
wire [0:104] sb_1__1__3_chany_top_out;
wire [0:0] sb_1__1__4_ccff_tail;
wire [0:104] sb_1__1__4_chanx_left_out;
wire [0:104] sb_1__1__4_chanx_right_out;
wire [0:104] sb_1__1__4_chany_bottom_out;
wire [0:104] sb_1__1__4_chany_top_out;
wire [0:0] sb_1__1__5_ccff_tail;
wire [0:104] sb_1__1__5_chanx_left_out;
wire [0:104] sb_1__1__5_chanx_right_out;
wire [0:104] sb_1__1__5_chany_bottom_out;
wire [0:104] sb_1__1__5_chany_top_out;
wire [0:0] sb_1__1__6_ccff_tail;
wire [0:104] sb_1__1__6_chanx_left_out;
wire [0:104] sb_1__1__6_chanx_right_out;
wire [0:104] sb_1__1__6_chany_bottom_out;
wire [0:104] sb_1__1__6_chany_top_out;
wire [0:0] sb_1__1__7_ccff_tail;
wire [0:104] sb_1__1__7_chanx_left_out;
wire [0:104] sb_1__1__7_chanx_right_out;
wire [0:104] sb_1__1__7_chany_bottom_out;
wire [0:104] sb_1__1__7_chany_top_out;
wire [0:0] sb_1__1__8_ccff_tail;
wire [0:104] sb_1__1__8_chanx_left_out;
wire [0:104] sb_1__1__8_chanx_right_out;
wire [0:104] sb_1__1__8_chany_bottom_out;
wire [0:104] sb_1__1__8_chany_top_out;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:104] sb_1__2__0_chanx_left_out;
wire [0:104] sb_1__2__0_chanx_right_out;
wire [0:104] sb_1__2__0_chany_bottom_out;
wire [0:104] sb_1__2__0_chany_top_out;
wire [0:0] sb_1__2__1_ccff_tail;
wire [0:104] sb_1__2__1_chanx_left_out;
wire [0:104] sb_1__2__1_chanx_right_out;
wire [0:104] sb_1__2__1_chany_bottom_out;
wire [0:104] sb_1__2__1_chany_top_out;
wire [0:0] sb_1__2__2_ccff_tail;
wire [0:104] sb_1__2__2_chanx_left_out;
wire [0:104] sb_1__2__2_chanx_right_out;
wire [0:104] sb_1__2__2_chany_bottom_out;
wire [0:104] sb_1__2__2_chany_top_out;
wire [0:0] sb_1__2__3_ccff_tail;
wire [0:104] sb_1__2__3_chanx_left_out;
wire [0:104] sb_1__2__3_chanx_right_out;
wire [0:104] sb_1__2__3_chany_bottom_out;
wire [0:104] sb_1__2__3_chany_top_out;
wire [0:0] sb_1__2__4_ccff_tail;
wire [0:104] sb_1__2__4_chanx_left_out;
wire [0:104] sb_1__2__4_chanx_right_out;
wire [0:104] sb_1__2__4_chany_bottom_out;
wire [0:104] sb_1__2__4_chany_top_out;
wire [0:0] sb_1__2__5_ccff_tail;
wire [0:104] sb_1__2__5_chanx_left_out;
wire [0:104] sb_1__2__5_chanx_right_out;
wire [0:104] sb_1__2__5_chany_bottom_out;
wire [0:104] sb_1__2__5_chany_top_out;
wire [0:0] sb_1__2__6_ccff_tail;
wire [0:104] sb_1__2__6_chanx_left_out;
wire [0:104] sb_1__2__6_chanx_right_out;
wire [0:104] sb_1__2__6_chany_bottom_out;
wire [0:104] sb_1__2__6_chany_top_out;
wire [0:0] sb_1__2__7_ccff_tail;
wire [0:104] sb_1__2__7_chanx_left_out;
wire [0:104] sb_1__2__7_chanx_right_out;
wire [0:104] sb_1__2__7_chany_bottom_out;
wire [0:104] sb_1__2__7_chany_top_out;
wire [0:0] sb_1__2__8_ccff_tail;
wire [0:104] sb_1__2__8_chanx_left_out;
wire [0:104] sb_1__2__8_chanx_right_out;
wire [0:104] sb_1__2__8_chany_bottom_out;
wire [0:104] sb_1__2__8_chany_top_out;
wire [0:0] sb_1__3__0_ccff_tail;
wire [0:104] sb_1__3__0_chanx_left_out;
wire [0:104] sb_1__3__0_chanx_right_out;
wire [0:104] sb_1__3__0_chany_bottom_out;
wire [0:104] sb_1__3__0_chany_top_out;
wire [0:0] sb_1__3__10_ccff_tail;
wire [0:104] sb_1__3__10_chanx_left_out;
wire [0:104] sb_1__3__10_chanx_right_out;
wire [0:104] sb_1__3__10_chany_bottom_out;
wire [0:104] sb_1__3__10_chany_top_out;
wire [0:0] sb_1__3__11_ccff_tail;
wire [0:104] sb_1__3__11_chanx_left_out;
wire [0:104] sb_1__3__11_chanx_right_out;
wire [0:104] sb_1__3__11_chany_bottom_out;
wire [0:104] sb_1__3__11_chany_top_out;
wire [0:0] sb_1__3__12_ccff_tail;
wire [0:104] sb_1__3__12_chanx_left_out;
wire [0:104] sb_1__3__12_chanx_right_out;
wire [0:104] sb_1__3__12_chany_bottom_out;
wire [0:104] sb_1__3__12_chany_top_out;
wire [0:0] sb_1__3__13_ccff_tail;
wire [0:104] sb_1__3__13_chanx_left_out;
wire [0:104] sb_1__3__13_chanx_right_out;
wire [0:104] sb_1__3__13_chany_bottom_out;
wire [0:104] sb_1__3__13_chany_top_out;
wire [0:0] sb_1__3__14_ccff_tail;
wire [0:104] sb_1__3__14_chanx_left_out;
wire [0:104] sb_1__3__14_chanx_right_out;
wire [0:104] sb_1__3__14_chany_bottom_out;
wire [0:104] sb_1__3__14_chany_top_out;
wire [0:0] sb_1__3__15_ccff_tail;
wire [0:104] sb_1__3__15_chanx_left_out;
wire [0:104] sb_1__3__15_chanx_right_out;
wire [0:104] sb_1__3__15_chany_bottom_out;
wire [0:104] sb_1__3__15_chany_top_out;
wire [0:0] sb_1__3__16_ccff_tail;
wire [0:104] sb_1__3__16_chanx_left_out;
wire [0:104] sb_1__3__16_chanx_right_out;
wire [0:104] sb_1__3__16_chany_bottom_out;
wire [0:104] sb_1__3__16_chany_top_out;
wire [0:0] sb_1__3__17_ccff_tail;
wire [0:104] sb_1__3__17_chanx_left_out;
wire [0:104] sb_1__3__17_chanx_right_out;
wire [0:104] sb_1__3__17_chany_bottom_out;
wire [0:104] sb_1__3__17_chany_top_out;
wire [0:0] sb_1__3__18_ccff_tail;
wire [0:104] sb_1__3__18_chanx_left_out;
wire [0:104] sb_1__3__18_chanx_right_out;
wire [0:104] sb_1__3__18_chany_bottom_out;
wire [0:104] sb_1__3__18_chany_top_out;
wire [0:0] sb_1__3__19_ccff_tail;
wire [0:104] sb_1__3__19_chanx_left_out;
wire [0:104] sb_1__3__19_chanx_right_out;
wire [0:104] sb_1__3__19_chany_bottom_out;
wire [0:104] sb_1__3__19_chany_top_out;
wire [0:0] sb_1__3__1_ccff_tail;
wire [0:104] sb_1__3__1_chanx_left_out;
wire [0:104] sb_1__3__1_chanx_right_out;
wire [0:104] sb_1__3__1_chany_bottom_out;
wire [0:104] sb_1__3__1_chany_top_out;
wire [0:0] sb_1__3__20_ccff_tail;
wire [0:104] sb_1__3__20_chanx_left_out;
wire [0:104] sb_1__3__20_chanx_right_out;
wire [0:104] sb_1__3__20_chany_bottom_out;
wire [0:104] sb_1__3__20_chany_top_out;
wire [0:0] sb_1__3__21_ccff_tail;
wire [0:104] sb_1__3__21_chanx_left_out;
wire [0:104] sb_1__3__21_chanx_right_out;
wire [0:104] sb_1__3__21_chany_bottom_out;
wire [0:104] sb_1__3__21_chany_top_out;
wire [0:0] sb_1__3__22_ccff_tail;
wire [0:104] sb_1__3__22_chanx_left_out;
wire [0:104] sb_1__3__22_chanx_right_out;
wire [0:104] sb_1__3__22_chany_bottom_out;
wire [0:104] sb_1__3__22_chany_top_out;
wire [0:0] sb_1__3__23_ccff_tail;
wire [0:104] sb_1__3__23_chanx_left_out;
wire [0:104] sb_1__3__23_chanx_right_out;
wire [0:104] sb_1__3__23_chany_bottom_out;
wire [0:104] sb_1__3__23_chany_top_out;
wire [0:0] sb_1__3__24_ccff_tail;
wire [0:104] sb_1__3__24_chanx_left_out;
wire [0:104] sb_1__3__24_chanx_right_out;
wire [0:104] sb_1__3__24_chany_bottom_out;
wire [0:104] sb_1__3__24_chany_top_out;
wire [0:0] sb_1__3__25_ccff_tail;
wire [0:104] sb_1__3__25_chanx_left_out;
wire [0:104] sb_1__3__25_chanx_right_out;
wire [0:104] sb_1__3__25_chany_bottom_out;
wire [0:104] sb_1__3__25_chany_top_out;
wire [0:0] sb_1__3__26_ccff_tail;
wire [0:104] sb_1__3__26_chanx_left_out;
wire [0:104] sb_1__3__26_chanx_right_out;
wire [0:104] sb_1__3__26_chany_bottom_out;
wire [0:104] sb_1__3__26_chany_top_out;
wire [0:0] sb_1__3__27_ccff_tail;
wire [0:104] sb_1__3__27_chanx_left_out;
wire [0:104] sb_1__3__27_chanx_right_out;
wire [0:104] sb_1__3__27_chany_bottom_out;
wire [0:104] sb_1__3__27_chany_top_out;
wire [0:0] sb_1__3__28_ccff_tail;
wire [0:104] sb_1__3__28_chanx_left_out;
wire [0:104] sb_1__3__28_chanx_right_out;
wire [0:104] sb_1__3__28_chany_bottom_out;
wire [0:104] sb_1__3__28_chany_top_out;
wire [0:0] sb_1__3__29_ccff_tail;
wire [0:104] sb_1__3__29_chanx_left_out;
wire [0:104] sb_1__3__29_chanx_right_out;
wire [0:104] sb_1__3__29_chany_bottom_out;
wire [0:104] sb_1__3__29_chany_top_out;
wire [0:0] sb_1__3__2_ccff_tail;
wire [0:104] sb_1__3__2_chanx_left_out;
wire [0:104] sb_1__3__2_chanx_right_out;
wire [0:104] sb_1__3__2_chany_bottom_out;
wire [0:104] sb_1__3__2_chany_top_out;
wire [0:0] sb_1__3__30_ccff_tail;
wire [0:104] sb_1__3__30_chanx_left_out;
wire [0:104] sb_1__3__30_chanx_right_out;
wire [0:104] sb_1__3__30_chany_bottom_out;
wire [0:104] sb_1__3__30_chany_top_out;
wire [0:0] sb_1__3__31_ccff_tail;
wire [0:104] sb_1__3__31_chanx_left_out;
wire [0:104] sb_1__3__31_chanx_right_out;
wire [0:104] sb_1__3__31_chany_bottom_out;
wire [0:104] sb_1__3__31_chany_top_out;
wire [0:0] sb_1__3__32_ccff_tail;
wire [0:104] sb_1__3__32_chanx_left_out;
wire [0:104] sb_1__3__32_chanx_right_out;
wire [0:104] sb_1__3__32_chany_bottom_out;
wire [0:104] sb_1__3__32_chany_top_out;
wire [0:0] sb_1__3__33_ccff_tail;
wire [0:104] sb_1__3__33_chanx_left_out;
wire [0:104] sb_1__3__33_chanx_right_out;
wire [0:104] sb_1__3__33_chany_bottom_out;
wire [0:104] sb_1__3__33_chany_top_out;
wire [0:0] sb_1__3__34_ccff_tail;
wire [0:104] sb_1__3__34_chanx_left_out;
wire [0:104] sb_1__3__34_chanx_right_out;
wire [0:104] sb_1__3__34_chany_bottom_out;
wire [0:104] sb_1__3__34_chany_top_out;
wire [0:0] sb_1__3__35_ccff_tail;
wire [0:104] sb_1__3__35_chanx_left_out;
wire [0:104] sb_1__3__35_chanx_right_out;
wire [0:104] sb_1__3__35_chany_bottom_out;
wire [0:104] sb_1__3__35_chany_top_out;
wire [0:0] sb_1__3__36_ccff_tail;
wire [0:104] sb_1__3__36_chanx_left_out;
wire [0:104] sb_1__3__36_chanx_right_out;
wire [0:104] sb_1__3__36_chany_bottom_out;
wire [0:104] sb_1__3__36_chany_top_out;
wire [0:0] sb_1__3__37_ccff_tail;
wire [0:104] sb_1__3__37_chanx_left_out;
wire [0:104] sb_1__3__37_chanx_right_out;
wire [0:104] sb_1__3__37_chany_bottom_out;
wire [0:104] sb_1__3__37_chany_top_out;
wire [0:0] sb_1__3__38_ccff_tail;
wire [0:104] sb_1__3__38_chanx_left_out;
wire [0:104] sb_1__3__38_chanx_right_out;
wire [0:104] sb_1__3__38_chany_bottom_out;
wire [0:104] sb_1__3__38_chany_top_out;
wire [0:0] sb_1__3__39_ccff_tail;
wire [0:104] sb_1__3__39_chanx_left_out;
wire [0:104] sb_1__3__39_chanx_right_out;
wire [0:104] sb_1__3__39_chany_bottom_out;
wire [0:104] sb_1__3__39_chany_top_out;
wire [0:0] sb_1__3__3_ccff_tail;
wire [0:104] sb_1__3__3_chanx_left_out;
wire [0:104] sb_1__3__3_chanx_right_out;
wire [0:104] sb_1__3__3_chany_bottom_out;
wire [0:104] sb_1__3__3_chany_top_out;
wire [0:0] sb_1__3__40_ccff_tail;
wire [0:104] sb_1__3__40_chanx_left_out;
wire [0:104] sb_1__3__40_chanx_right_out;
wire [0:104] sb_1__3__40_chany_bottom_out;
wire [0:104] sb_1__3__40_chany_top_out;
wire [0:0] sb_1__3__41_ccff_tail;
wire [0:104] sb_1__3__41_chanx_left_out;
wire [0:104] sb_1__3__41_chanx_right_out;
wire [0:104] sb_1__3__41_chany_bottom_out;
wire [0:104] sb_1__3__41_chany_top_out;
wire [0:0] sb_1__3__42_ccff_tail;
wire [0:104] sb_1__3__42_chanx_left_out;
wire [0:104] sb_1__3__42_chanx_right_out;
wire [0:104] sb_1__3__42_chany_bottom_out;
wire [0:104] sb_1__3__42_chany_top_out;
wire [0:0] sb_1__3__43_ccff_tail;
wire [0:104] sb_1__3__43_chanx_left_out;
wire [0:104] sb_1__3__43_chanx_right_out;
wire [0:104] sb_1__3__43_chany_bottom_out;
wire [0:104] sb_1__3__43_chany_top_out;
wire [0:0] sb_1__3__44_ccff_tail;
wire [0:104] sb_1__3__44_chanx_left_out;
wire [0:104] sb_1__3__44_chanx_right_out;
wire [0:104] sb_1__3__44_chany_bottom_out;
wire [0:104] sb_1__3__44_chany_top_out;
wire [0:0] sb_1__3__45_ccff_tail;
wire [0:104] sb_1__3__45_chanx_left_out;
wire [0:104] sb_1__3__45_chanx_right_out;
wire [0:104] sb_1__3__45_chany_bottom_out;
wire [0:104] sb_1__3__45_chany_top_out;
wire [0:0] sb_1__3__46_ccff_tail;
wire [0:104] sb_1__3__46_chanx_left_out;
wire [0:104] sb_1__3__46_chanx_right_out;
wire [0:104] sb_1__3__46_chany_bottom_out;
wire [0:104] sb_1__3__46_chany_top_out;
wire [0:0] sb_1__3__47_ccff_tail;
wire [0:104] sb_1__3__47_chanx_left_out;
wire [0:104] sb_1__3__47_chanx_right_out;
wire [0:104] sb_1__3__47_chany_bottom_out;
wire [0:104] sb_1__3__47_chany_top_out;
wire [0:0] sb_1__3__48_ccff_tail;
wire [0:104] sb_1__3__48_chanx_left_out;
wire [0:104] sb_1__3__48_chanx_right_out;
wire [0:104] sb_1__3__48_chany_bottom_out;
wire [0:104] sb_1__3__48_chany_top_out;
wire [0:0] sb_1__3__49_ccff_tail;
wire [0:104] sb_1__3__49_chanx_left_out;
wire [0:104] sb_1__3__49_chanx_right_out;
wire [0:104] sb_1__3__49_chany_bottom_out;
wire [0:104] sb_1__3__49_chany_top_out;
wire [0:0] sb_1__3__4_ccff_tail;
wire [0:104] sb_1__3__4_chanx_left_out;
wire [0:104] sb_1__3__4_chanx_right_out;
wire [0:104] sb_1__3__4_chany_bottom_out;
wire [0:104] sb_1__3__4_chany_top_out;
wire [0:0] sb_1__3__50_ccff_tail;
wire [0:104] sb_1__3__50_chanx_left_out;
wire [0:104] sb_1__3__50_chanx_right_out;
wire [0:104] sb_1__3__50_chany_bottom_out;
wire [0:104] sb_1__3__50_chany_top_out;
wire [0:0] sb_1__3__51_ccff_tail;
wire [0:104] sb_1__3__51_chanx_left_out;
wire [0:104] sb_1__3__51_chanx_right_out;
wire [0:104] sb_1__3__51_chany_bottom_out;
wire [0:104] sb_1__3__51_chany_top_out;
wire [0:0] sb_1__3__52_ccff_tail;
wire [0:104] sb_1__3__52_chanx_left_out;
wire [0:104] sb_1__3__52_chanx_right_out;
wire [0:104] sb_1__3__52_chany_bottom_out;
wire [0:104] sb_1__3__52_chany_top_out;
wire [0:0] sb_1__3__53_ccff_tail;
wire [0:104] sb_1__3__53_chanx_left_out;
wire [0:104] sb_1__3__53_chanx_right_out;
wire [0:104] sb_1__3__53_chany_bottom_out;
wire [0:104] sb_1__3__53_chany_top_out;
wire [0:0] sb_1__3__54_ccff_tail;
wire [0:104] sb_1__3__54_chanx_left_out;
wire [0:104] sb_1__3__54_chanx_right_out;
wire [0:104] sb_1__3__54_chany_bottom_out;
wire [0:104] sb_1__3__54_chany_top_out;
wire [0:0] sb_1__3__55_ccff_tail;
wire [0:104] sb_1__3__55_chanx_left_out;
wire [0:104] sb_1__3__55_chanx_right_out;
wire [0:104] sb_1__3__55_chany_bottom_out;
wire [0:104] sb_1__3__55_chany_top_out;
wire [0:0] sb_1__3__56_ccff_tail;
wire [0:104] sb_1__3__56_chanx_left_out;
wire [0:104] sb_1__3__56_chanx_right_out;
wire [0:104] sb_1__3__56_chany_bottom_out;
wire [0:104] sb_1__3__56_chany_top_out;
wire [0:0] sb_1__3__5_ccff_tail;
wire [0:104] sb_1__3__5_chanx_left_out;
wire [0:104] sb_1__3__5_chanx_right_out;
wire [0:104] sb_1__3__5_chany_bottom_out;
wire [0:104] sb_1__3__5_chany_top_out;
wire [0:0] sb_1__3__6_ccff_tail;
wire [0:104] sb_1__3__6_chanx_left_out;
wire [0:104] sb_1__3__6_chanx_right_out;
wire [0:104] sb_1__3__6_chany_bottom_out;
wire [0:104] sb_1__3__6_chany_top_out;
wire [0:0] sb_1__3__7_ccff_tail;
wire [0:104] sb_1__3__7_chanx_left_out;
wire [0:104] sb_1__3__7_chanx_right_out;
wire [0:104] sb_1__3__7_chany_bottom_out;
wire [0:104] sb_1__3__7_chany_top_out;
wire [0:0] sb_1__3__8_ccff_tail;
wire [0:104] sb_1__3__8_chanx_left_out;
wire [0:104] sb_1__3__8_chanx_right_out;
wire [0:104] sb_1__3__8_chany_bottom_out;
wire [0:104] sb_1__3__8_chany_top_out;
wire [0:0] sb_1__3__9_ccff_tail;
wire [0:104] sb_1__3__9_chanx_left_out;
wire [0:104] sb_1__3__9_chanx_right_out;
wire [0:104] sb_1__3__9_chany_bottom_out;
wire [0:104] sb_1__3__9_chany_top_out;
wire [0:0] sb_5__5__0_ccff_tail;
wire [0:104] sb_5__5__0_chanx_left_out;
wire [0:104] sb_5__5__0_chanx_right_out;
wire [0:104] sb_5__5__0_chany_bottom_out;
wire [0:104] sb_5__5__0_chany_top_out;
wire [0:0] sb_5__5__1_ccff_tail;
wire [0:104] sb_5__5__1_chanx_left_out;
wire [0:104] sb_5__5__1_chanx_right_out;
wire [0:104] sb_5__5__1_chany_bottom_out;
wire [0:104] sb_5__5__1_chany_top_out;
wire [0:0] sb_5__6__0_ccff_tail;
wire [0:104] sb_5__6__0_chanx_left_out;
wire [0:104] sb_5__6__0_chanx_right_out;
wire [0:104] sb_5__6__0_chany_bottom_out;
wire [0:104] sb_5__6__0_chany_top_out;
wire [0:0] sb_5__6__1_ccff_tail;
wire [0:104] sb_5__6__1_chanx_left_out;
wire [0:104] sb_5__6__1_chanx_right_out;
wire [0:104] sb_5__6__1_chany_bottom_out;
wire [0:104] sb_5__6__1_chany_top_out;
wire [0:0] sb_6__5__0_ccff_tail;
wire [0:104] sb_6__5__0_chanx_left_out;
wire [0:104] sb_6__5__0_chanx_right_out;
wire [0:104] sb_6__5__0_chany_bottom_out;
wire [0:104] sb_6__5__0_chany_top_out;
wire [0:0] sb_6__6__0_ccff_tail;
wire [0:104] sb_6__6__0_chanx_left_out;
wire [0:104] sb_6__6__0_chanx_right_out;
wire [0:104] sb_6__6__0_chany_bottom_out;
wire [0:104] sb_6__6__0_chany_top_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_4__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_top grid_io_top_5__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_4_ccff_tail));

	grid_io_top grid_io_top_6__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_5_ccff_tail));

	grid_io_top grid_io_top_7__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__6_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_6_ccff_tail));

	grid_io_top grid_io_top_8__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__7_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_7_ccff_tail));

	grid_io_top grid_io_top_9__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__8_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_8_ccff_tail));

	grid_io_top grid_io_top_10__11_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__10__9_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_9_ccff_tail));

	grid_io_right grid_io_right_11__10_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_11__9_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_11__8_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_11__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right grid_io_right_11__6_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right grid_io_right_11__5_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_right grid_io_right_11__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[128:135]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_6_ccff_tail));

	grid_io_right grid_io_right_11__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[136:143]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_8_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_7_ccff_tail));

	grid_io_right grid_io_right_11__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[144:151]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_9_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_8_ccff_tail));

	grid_io_right grid_io_right_11__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[152:159]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_9_ccff_tail));

	grid_io_bottom grid_io_bottom_10__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[160:167]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_9__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[168:175]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_8__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[176:183]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_7__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[184:191]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_bottom grid_io_bottom_6__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[192:199]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_4_ccff_tail));

	grid_io_bottom grid_io_bottom_5__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[200:207]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_5_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[208:215]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_6_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[216:223]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_7_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[224:231]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_8_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[232:239]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_9_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[240:247]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[248:255]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[256:263]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[264:271]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[272:279]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[280:287]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_io_left grid_io_left_0__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[288:295]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_6_ccff_tail));

	grid_io_left grid_io_left_0__8_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[296:303]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_7_ccff_tail));

	grid_io_left grid_io_left_0__9_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[304:311]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_8_ccff_tail));

	grid_io_left grid_io_left_0__10_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[312:319]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__3__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_9_ccff_tail));

	grid_io grid_io_1__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[320:327]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_0_ccff_tail));

	grid_io grid_io_1__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[328:335]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_1_ccff_tail));

	grid_io grid_io_2__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[408:415]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_2_ccff_tail));

	grid_io grid_io_2__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[416:423]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_3_ccff_tail));

	grid_io grid_io_3__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[400:407]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_4_ccff_tail));

	grid_io grid_io_3__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[472:479]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_5_ccff_tail));

	grid_io grid_io_4__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[392:399]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_6_ccff_tail));

	grid_io grid_io_4__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[464:471]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_7_ccff_tail));

	grid_io grid_io_5__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[384:391]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_8_ccff_tail));

	grid_io grid_io_5__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[456:463]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_9_ccff_tail));

	grid_io grid_io_6__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[376:383]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_10_ccff_tail));

	grid_io grid_io_6__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[448:455]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_11_ccff_tail));

	grid_io grid_io_7__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[368:375]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_12_ccff_tail));

	grid_io grid_io_7__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[440:447]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_13_ccff_tail));

	grid_io grid_io_8__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[360:367]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_14_ccff_tail));

	grid_io grid_io_8__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[432:439]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_15_ccff_tail));

	grid_io grid_io_9__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[352:359]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_16_ccff_tail));

	grid_io grid_io_9__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[424:431]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_17_ccff_tail));

	grid_io grid_io_10__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[344:351]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_18_ccff_tail));

	grid_io grid_io_10__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[336:343]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_19_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_1__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_1__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_1__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_1__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_2__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_2__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_2__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_2__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_2__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_3__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_3__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_3__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__22_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_3__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__23_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__24_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_24_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__25_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_25_ccff_tail));

	grid_clb grid_clb_4__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__26_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_26_ccff_tail));

	grid_clb grid_clb_4__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__27_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_27_ccff_tail));

	grid_clb grid_clb_4__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__28_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_28_ccff_tail));

	grid_clb grid_clb_4__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__29_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_29_ccff_tail));

	grid_clb grid_clb_4__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__30_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_30_ccff_tail));

	grid_clb grid_clb_4__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__31_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_31_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__32_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_32_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__33_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_33_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__34_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_34_ccff_tail));

	grid_clb grid_clb_5__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_5__6__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_35_ccff_tail));

	grid_clb grid_clb_5__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__35_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_36_ccff_tail));

	grid_clb grid_clb_5__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__36_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_37_ccff_tail));

	grid_clb grid_clb_5__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__37_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_38_ccff_tail));

	grid_clb grid_clb_5__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_5__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__38_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_39_ccff_tail));

	grid_clb grid_clb_6__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__39_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_40_ccff_tail));

	grid_clb grid_clb_6__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__40_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_41_ccff_tail));

	grid_clb grid_clb_6__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__41_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_42_ccff_tail));

	grid_clb grid_clb_6__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__42_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_43_ccff_tail));

	grid_clb grid_clb_6__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__43_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_44_ccff_tail));

	grid_clb grid_clb_6__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__44_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_45_ccff_tail));

	grid_clb grid_clb_6__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_6__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__45_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_46_ccff_tail));

	grid_clb grid_clb_7__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__46_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_47_ccff_tail));

	grid_clb grid_clb_7__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__47_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_48_ccff_tail));

	grid_clb grid_clb_7__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__48_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_49_ccff_tail));

	grid_clb grid_clb_7__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__49_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_50_ccff_tail));

	grid_clb grid_clb_7__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__50_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_51_ccff_tail));

	grid_clb grid_clb_7__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__51_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_52_ccff_tail));

	grid_clb grid_clb_7__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__52_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_53_ccff_tail));

	grid_clb grid_clb_7__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_7__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__53_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_54_ccff_tail));

	grid_clb grid_clb_8__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__54_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_55_ccff_tail));

	grid_clb grid_clb_8__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__55_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_56_ccff_tail));

	grid_clb grid_clb_8__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__56_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_57_ccff_tail));

	grid_clb grid_clb_8__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__57_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_58_ccff_tail));

	grid_clb grid_clb_8__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__58_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_59_ccff_tail));

	grid_clb grid_clb_8__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__59_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_60_ccff_tail));

	grid_clb grid_clb_8__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__60_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_61_ccff_tail));

	grid_clb grid_clb_8__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_8__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__61_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_62_ccff_tail));

	grid_clb grid_clb_9__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__62_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_63_ccff_tail));

	grid_clb grid_clb_9__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__63_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_64_ccff_tail));

	grid_clb grid_clb_9__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__64_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_65_ccff_tail));

	grid_clb grid_clb_9__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_5__6__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_66_ccff_tail));

	grid_clb grid_clb_9__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__65_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_67_ccff_tail));

	grid_clb grid_clb_9__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__66_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_68_ccff_tail));

	grid_clb grid_clb_9__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__67_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_69_ccff_tail));

	grid_clb grid_clb_9__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_9__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__3__68_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_70_ccff_tail));

	grid_clb grid_clb_10__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_71_ccff_tail));

	grid_clb grid_clb_10__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_72_ccff_tail));

	grid_clb grid_clb_10__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_73_ccff_tail));

	grid_clb grid_clb_10__7_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__7__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_74_ccff_tail));

	grid_clb grid_clb_10__8_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__8__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_75_ccff_tail));

	grid_clb grid_clb_10__9_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__9__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_76_ccff_tail));

	grid_clb grid_clb_10__10_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_10__10__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_10__3__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_77_ccff_tail));

	grid_router grid_router_6__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_6__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	grid_router grid_router_10__6_ (
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_rst__0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.right_width_0_height_0_subtile_0__pin_clk_0_(grid_router_10__6__undriven_right_width_0_height_0_subtile_0__pin_clk_0_),
		.bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:104]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:104]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:104]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__2_ sb_0__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__2__0_chany_top_out[0:104]),
		.chanx_right_out(sb_0__2__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__2__0_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__2__0_ccff_tail));

	sb_0__3_ sb_0__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__1_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_0__3__0_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__0_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__0_ccff_tail));

	sb_0__3_ sb_0__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__2_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__1_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_0__3__1_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__1_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__1_ccff_tail));

	sb_0__3_ sb_0__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__3_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__2_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__2_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_6_ccff_tail),
		.chany_top_out(sb_0__3__2_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__2_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__2_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__2_ccff_tail));

	sb_0__3_ sb_0__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__4_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__3_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__3_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_7_ccff_tail),
		.chany_top_out(sb_0__3__3_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__3_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__3_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__3_ccff_tail));

	sb_0__3_ sb_0__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__5_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__4_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__4_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_8_ccff_tail),
		.chany_top_out(sb_0__3__4_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__4_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__4_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__4_ccff_tail));

	sb_0__3_ sb_0__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__6_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__5_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__5_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_9_ccff_tail),
		.chany_top_out(sb_0__3__5_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__5_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__5_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__5_ccff_tail));

	sb_0__3_ sb_0__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__3__7_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__6_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__6_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__10__0_ccff_tail),
		.chany_top_out(sb_0__3__6_chany_top_out[0:104]),
		.chanx_right_out(sb_0__3__6_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__3__6_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__3__6_ccff_tail));

	sb_0__10_ sb_0__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__3__7_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__10__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_0__10__0_chany_bottom_out[0:104]),
		.ccff_tail(sb_0__10__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_2_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__8_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__8_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_4_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_5__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__10_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__10_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__8_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_6_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__0_ sb_6__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__12_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__12_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__10_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_8_ccff_tail),
		.chany_top_out(sb_1__0__5_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__5_ccff_tail));

	sb_1__0_ sb_7__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__14_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__14_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__12_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_10_ccff_tail),
		.chany_top_out(sb_1__0__6_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__6_ccff_tail));

	sb_1__0_ sb_8__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__16_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__16_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__14_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_12_ccff_tail),
		.chany_top_out(sb_1__0__7_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__7_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__7_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__7_ccff_tail));

	sb_1__0_ sb_9__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__18_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__18_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__16_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_14_ccff_tail),
		.chany_top_out(sb_1__0__8_chany_top_out[0:104]),
		.chanx_right_out(sb_1__0__8_chanx_right_out[0:104]),
		.chanx_left_out(sb_1__0__8_chanx_left_out[0:104]),
		.ccff_tail(sb_1__0__8_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_3_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_5_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_4_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_7_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_4__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__9_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__9_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__8_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_6_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_9_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_5__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__11_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__11_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__10_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__9_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_8_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_11_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_6__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__13_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__13_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__12_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__11_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_10_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_13_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_7__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__15_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__15_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__14_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__13_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_12_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_15_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_8__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__17_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__17_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__16_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__15_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_14_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_17_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_9__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__19_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__19_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__18_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__17_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_16_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_19_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:104]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:104]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_1_ccff_tail),
		.chany_top_out(sb_1__2__0_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_1__2_ sb_2__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__8_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__2_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__2__1_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__1_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__1_ccff_tail));

	sb_1__2_ sb_3__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__16_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__3_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__2_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_5_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__2__2_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__2_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__2_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__2_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__2_ccff_tail));

	sb_1__2_ sb_4__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__24_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__4_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__9_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__3_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_7_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__2__3_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__3_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__3_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__3_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__3_ccff_tail));

	sb_1__2_ sb_5__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__32_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__5_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__11_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__4_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_9_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_24_ccff_tail),
		.chany_top_out(sb_1__2__4_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__4_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__4_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__4_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__4_ccff_tail));

	sb_1__2_ sb_6__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__39_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__6_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__13_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__5_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_11_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_32_ccff_tail),
		.chany_top_out(sb_1__2__5_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__5_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__5_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__5_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__5_ccff_tail));

	sb_1__2_ sb_7__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__46_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__7_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__15_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__6_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_13_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_40_ccff_tail),
		.chany_top_out(sb_1__2__6_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__6_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__6_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__6_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__6_ccff_tail));

	sb_1__2_ sb_8__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__54_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__8_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__17_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__7_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_15_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_47_ccff_tail),
		.chany_top_out(sb_1__2__7_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__7_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__7_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__7_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__7_ccff_tail));

	sb_1__2_ sb_9__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__62_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__9_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__19_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__8_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_17_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_55_ccff_tail),
		.chany_top_out(sb_1__2__8_chany_top_out[0:104]),
		.chanx_right_out(sb_1__2__8_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__2__8_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__2__8_chanx_left_out[0:104]),
		.ccff_tail(sb_1__2__8_ccff_tail));

	sb_1__3_ sb_1__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__1_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__7_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__3__0_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__0_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__0_ccff_tail));

	sb_1__3_ sb_1__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__2_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__8_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__1_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__3__1_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__1_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__1_ccff_tail));

	sb_1__3_ sb_1__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__3_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__9_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__2_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__2_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__3__2_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__2_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__2_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__2_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__2_ccff_tail));

	sb_1__3_ sb_1__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__4_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__10_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__3_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__3_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__3__3_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__3_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__3_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__3_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__3_ccff_tail));

	sb_1__3_ sb_1__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__5_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__11_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__4_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__4_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__3__4_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__4_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__4_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__4_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__4_ccff_tail));

	sb_1__3_ sb_1__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__6_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__12_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__5_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__5_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__3__5_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__5_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__5_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__5_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__5_ccff_tail));

	sb_1__3_ sb_1__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__7_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__13_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__6_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__6_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__3__6_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__6_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__6_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__6_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__6_ccff_tail));

	sb_1__3_ sb_2__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__9_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__14_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__8_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__7_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_1__3__7_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__7_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__7_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__7_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__7_ccff_tail));

	sb_1__3_ sb_2__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__10_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__15_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__9_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__8_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__3__8_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__8_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__8_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__8_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__8_ccff_tail));

	sb_1__3_ sb_2__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__11_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__16_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__10_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__9_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_1__3__9_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__9_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__9_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__9_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__9_ccff_tail));

	sb_1__3_ sb_2__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__12_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__17_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__11_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__10_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__3__10_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__10_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__10_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__10_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__10_ccff_tail));

	sb_1__3_ sb_2__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__13_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__18_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__12_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__11_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_1__3__11_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__11_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__11_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__11_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__11_ccff_tail));

	sb_1__3_ sb_2__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__14_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__19_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__13_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__12_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__3__12_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__12_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__12_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__12_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__12_ccff_tail));

	sb_1__3_ sb_2__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__15_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__20_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__14_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__13_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_1__3__13_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__13_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__13_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__13_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__13_ccff_tail));

	sb_1__3_ sb_3__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__17_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__21_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__16_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__14_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_25_ccff_tail),
		.chany_top_out(sb_1__3__14_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__14_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__14_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__14_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__14_ccff_tail));

	sb_1__3_ sb_3__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__18_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__22_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__17_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__15_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__3__15_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__15_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__15_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__15_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__15_ccff_tail));

	sb_1__3_ sb_3__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__19_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__23_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__18_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__16_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_27_ccff_tail),
		.chany_top_out(sb_1__3__16_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__16_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__16_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__16_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__16_ccff_tail));

	sb_1__3_ sb_3__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__20_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__24_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__19_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__17_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__3__17_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__17_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__17_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__17_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__17_ccff_tail));

	sb_1__3_ sb_3__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__21_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__25_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__20_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__18_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_29_ccff_tail),
		.chany_top_out(sb_1__3__18_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__18_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__18_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__18_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__18_ccff_tail));

	sb_1__3_ sb_3__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__22_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__26_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__21_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__19_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__3__19_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__19_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__19_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__19_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__19_ccff_tail));

	sb_1__3_ sb_3__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__23_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__27_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__22_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__20_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_31_ccff_tail),
		.chany_top_out(sb_1__3__20_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__20_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__20_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__20_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__20_ccff_tail));

	sb_1__3_ sb_4__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__25_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__28_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__24_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__21_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_33_ccff_tail),
		.chany_top_out(sb_1__3__21_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__21_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__21_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__21_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__21_ccff_tail));

	sb_1__3_ sb_4__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__26_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__29_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__25_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__22_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__3__22_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__22_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__22_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__22_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__22_ccff_tail));

	sb_1__3_ sb_4__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__27_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__30_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__26_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__23_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_35_ccff_tail),
		.chany_top_out(sb_1__3__23_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__23_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__23_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__23_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__23_ccff_tail));

	sb_1__3_ sb_4__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__28_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__31_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__27_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__24_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_1__3__24_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__24_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__24_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__24_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__24_ccff_tail));

	sb_1__3_ sb_4__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__29_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__32_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__28_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__25_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_37_ccff_tail),
		.chany_top_out(sb_1__3__25_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__25_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__25_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__25_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__25_ccff_tail));

	sb_1__3_ sb_4__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__30_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__33_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__29_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__26_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_1__3__26_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__26_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__26_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__26_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__26_ccff_tail));

	sb_1__3_ sb_4__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__31_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__34_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__30_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__27_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_39_ccff_tail),
		.chany_top_out(sb_1__3__27_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__27_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__27_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__27_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__27_ccff_tail));

	sb_1__3_ sb_5__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__33_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__35_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__32_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__28_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_41_ccff_tail),
		.chany_top_out(sb_1__3__28_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__28_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__28_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__28_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__28_ccff_tail));

	sb_1__3_ sb_5__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__34_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__36_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__33_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__29_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_26_ccff_tail),
		.chany_top_out(sb_1__3__29_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__29_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__29_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__29_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__29_ccff_tail));

	sb_1__3_ sb_5__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__36_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__37_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__35_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__32_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_44_ccff_tail),
		.chany_top_out(sb_1__3__30_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__30_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__30_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__30_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__30_ccff_tail));

	sb_1__3_ sb_5__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__37_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__38_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__36_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__33_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_30_ccff_tail),
		.chany_top_out(sb_1__3__31_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__31_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__31_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__31_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__31_ccff_tail));

	sb_1__3_ sb_5__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__38_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__39_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__37_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__34_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_46_ccff_tail),
		.chany_top_out(sb_1__3__32_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__32_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__32_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__32_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__32_ccff_tail));

	sb_1__3_ sb_6__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__40_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__40_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__39_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__35_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_48_ccff_tail),
		.chany_top_out(sb_1__3__33_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__33_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__33_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__33_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__33_ccff_tail));

	sb_1__3_ sb_6__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__41_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__41_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__40_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__36_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_34_ccff_tail),
		.chany_top_out(sb_1__3__34_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__34_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__34_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__34_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__34_ccff_tail));

	sb_1__3_ sb_6__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__43_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__44_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__42_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__37_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_52_ccff_tail),
		.chany_top_out(sb_1__3__35_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__35_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__35_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__35_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__35_ccff_tail));

	sb_1__3_ sb_6__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__44_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__45_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__43_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__38_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_38_ccff_tail),
		.chany_top_out(sb_1__3__36_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__36_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__36_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__36_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__36_ccff_tail));

	sb_1__3_ sb_6__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__45_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__46_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__44_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__39_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_54_ccff_tail),
		.chany_top_out(sb_1__3__37_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__37_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__37_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__37_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__37_ccff_tail));

	sb_1__3_ sb_7__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__47_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__47_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__46_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__40_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_56_ccff_tail),
		.chany_top_out(sb_1__3__38_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__38_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__38_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__38_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__38_ccff_tail));

	sb_1__3_ sb_7__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__48_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__48_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__47_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__41_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_42_ccff_tail),
		.chany_top_out(sb_1__3__39_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__39_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__39_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__39_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__39_ccff_tail));

	sb_1__3_ sb_7__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__49_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__49_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__48_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__42_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_58_ccff_tail),
		.chany_top_out(sb_1__3__40_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__40_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__40_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__40_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__40_ccff_tail));

	sb_1__3_ sb_7__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__50_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__50_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__49_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__43_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_43_ccff_tail),
		.chany_top_out(sb_1__3__41_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__41_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__41_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__41_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__41_ccff_tail));

	sb_1__3_ sb_7__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__51_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__51_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__50_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__44_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_60_ccff_tail),
		.chany_top_out(sb_1__3__42_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__42_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__42_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__42_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__42_ccff_tail));

	sb_1__3_ sb_7__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__52_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__52_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__51_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__45_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_45_ccff_tail),
		.chany_top_out(sb_1__3__43_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__43_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__43_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__43_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__43_ccff_tail));

	sb_1__3_ sb_7__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__53_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__53_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__52_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__46_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_62_ccff_tail),
		.chany_top_out(sb_1__3__44_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__44_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__44_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__44_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__44_ccff_tail));

	sb_1__3_ sb_8__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__55_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__54_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__54_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__47_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_64_ccff_tail),
		.chany_top_out(sb_1__3__45_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__45_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__45_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__45_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__45_ccff_tail));

	sb_1__3_ sb_8__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__56_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__55_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__55_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_64_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__48_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_49_ccff_tail),
		.chany_top_out(sb_1__3__46_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__46_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__46_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__46_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__46_ccff_tail));

	sb_1__3_ sb_8__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__57_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__56_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__56_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_65_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__49_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_66_ccff_tail),
		.chany_top_out(sb_1__3__47_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__47_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__47_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__47_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__47_ccff_tail));

	sb_1__3_ sb_8__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__58_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__57_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__57_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_66_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__50_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_51_ccff_tail),
		.chany_top_out(sb_1__3__48_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__48_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__48_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__48_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__48_ccff_tail));

	sb_1__3_ sb_8__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__59_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__58_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__58_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_67_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__51_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_68_ccff_tail),
		.chany_top_out(sb_1__3__49_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__49_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__49_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__49_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__49_ccff_tail));

	sb_1__3_ sb_8__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__60_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__59_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__59_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_68_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__52_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_53_ccff_tail),
		.chany_top_out(sb_1__3__50_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__50_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__50_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__50_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__50_ccff_tail));

	sb_1__3_ sb_8__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__61_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__60_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__60_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_69_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__53_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_70_ccff_tail),
		.chany_top_out(sb_1__3__51_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__51_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__51_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__51_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__51_ccff_tail));

	sb_1__3_ sb_9__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__63_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__61_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__62_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_71_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__54_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_64_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_72_ccff_tail),
		.chany_top_out(sb_1__3__52_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__52_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__52_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__52_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__52_ccff_tail));

	sb_1__3_ sb_9__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__64_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__62_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__63_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_72_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_64_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__55_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_65_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_64_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_57_ccff_tail),
		.chany_top_out(sb_1__3__53_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__53_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__53_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__53_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__53_ccff_tail));

	sb_1__3_ sb_9__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__66_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__63_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__65_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__58_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_68_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_67_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_75_ccff_tail),
		.chany_top_out(sb_1__3__54_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__54_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__54_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__54_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__54_ccff_tail));

	sb_1__3_ sb_9__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__67_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__64_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__66_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_75_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_68_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__59_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_69_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_68_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_61_ccff_tail),
		.chany_top_out(sb_1__3__55_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__55_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__55_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__55_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__55_ccff_tail));

	sb_1__3_ sb_9__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__68_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__65_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__67_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_76_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_69_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__60_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_70_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_69_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_77_ccff_tail),
		.chany_top_out(sb_1__3__56_chany_top_out[0:104]),
		.chanx_right_out(sb_1__3__56_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__3__56_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__3__56_chanx_left_out[0:104]),
		.ccff_tail(sb_1__3__56_ccff_tail));

	sb_1__10_ sb_1__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__7_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__10__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__0_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__0_ccff_tail));

	sb_1__10_ sb_2__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__2_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__15_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__10__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__1_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__1_ccff_tail));

	sb_1__10_ sb_3__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__3_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__23_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__2_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chanx_right_out(sb_1__10__2_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__2_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__2_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__2_ccff_tail));

	sb_1__10_ sb_4__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__4_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__31_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__3_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_4_ccff_tail),
		.chanx_right_out(sb_1__10__3_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__3_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__3_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__3_ccff_tail));

	sb_1__10_ sb_5__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__5_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__38_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__4_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_4_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_5_ccff_tail),
		.chanx_right_out(sb_1__10__4_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__4_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__4_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__4_ccff_tail));

	sb_1__10_ sb_6__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__6_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__45_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__5_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_5_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_6_ccff_tail),
		.chanx_right_out(sb_1__10__5_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__5_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__5_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__5_ccff_tail));

	sb_1__10_ sb_7__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__7_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__53_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__6_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_6_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_7_ccff_tail),
		.chanx_right_out(sb_1__10__6_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__6_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__6_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__6_ccff_tail));

	sb_1__10_ sb_8__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__8_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__61_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_70_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__7_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_7_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_8_ccff_tail),
		.chanx_right_out(sb_1__10__7_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__7_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__7_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__7_ccff_tail));

	sb_1__10_ sb_9__10_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__10__9_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__68_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_77_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_70_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__8_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_8_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_70_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_9_ccff_tail),
		.chanx_right_out(sb_1__10__8_chanx_right_out[0:104]),
		.chany_bottom_out(sb_1__10__8_chany_bottom_out[0:104]),
		.chanx_left_out(sb_1__10__8_chanx_left_out[0:104]),
		.ccff_tail(sb_1__10__8_ccff_tail));

	sb_5__5_ sb_5__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__6__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_6__5__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__34_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__30_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(cby_6__6__0_ccff_tail),
		.chany_top_out(sb_5__5__0_chany_top_out[0:104]),
		.chanx_right_out(sb_5__5__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_5__5__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_5__5__0_chanx_left_out[0:104]),
		.ccff_tail(sb_5__5__0_ccff_tail));

	sb_5__5_ sb_9__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_5__6__1_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.chanx_right_in(cbx_6__5__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__64_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_73_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_65_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__56_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_66_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_65_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(cby_10__6__0_ccff_tail),
		.chany_top_out(sb_5__5__1_chany_top_out[0:104]),
		.chanx_right_out(sb_5__5__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_5__5__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_5__5__1_chanx_left_out[0:104]),
		.ccff_tail(sb_5__5__1_ccff_tail));

	sb_5__6_ sb_5__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__35_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_6__6__0_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_5__6__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_0_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__31_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_28_ccff_tail),
		.chany_top_out(sb_5__6__0_chany_top_out[0:104]),
		.chanx_right_out(sb_5__6__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_5__6__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_5__6__0_chanx_left_out[0:104]),
		.ccff_tail(sb_5__6__0_ccff_tail));

	sb_5__6_ sb_9__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__65_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_67_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_74_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_6__6__1_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.chany_bottom_in(cby_5__6__1_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_0_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_2_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_6_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_10_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_14_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_18_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_22_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_26_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_30_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_1_34_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_7_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_11_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_15_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_19_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_23_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_27_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_2_31_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_4_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_8_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_12_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_16_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_20_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_24_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_28_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_3_32_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_odata_4_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_oack_4_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_1_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_ordy_3_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_0_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_2_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_(grid_router_1_left_width_0_height_0_subtile_0__pin_olck_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_66_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__57_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_67_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_66_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_59_ccff_tail),
		.chany_top_out(sb_5__6__1_chany_top_out[0:104]),
		.chanx_right_out(sb_5__6__1_chanx_right_out[0:104]),
		.chany_bottom_out(sb_5__6__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_5__6__1_chanx_left_out[0:104]),
		.ccff_tail(sb_5__6__1_ccff_tail));

	sb_6__5_ sb_6__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_6__6__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__42_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__3__41_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_6__5__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_50_ccff_tail),
		.chany_top_out(sb_6__5__0_chany_top_out[0:104]),
		.chanx_right_out(sb_6__5__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_6__5__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_6__5__0_chanx_left_out[0:104]),
		.ccff_tail(sb_6__5__0_ccff_tail));

	sb_6__6_ sb_6__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__3__42_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__43_chanx_left_out[0:104]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_6__6__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_6__6__0_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_0_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_0_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(grid_clb_36_ccff_tail),
		.chany_top_out(sb_6__6__0_chany_top_out[0:104]),
		.chanx_right_out(sb_6__6__0_chanx_right_out[0:104]),
		.chany_bottom_out(sb_6__6__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_6__6__0_chanx_left_out[0:104]),
		.ccff_tail(sb_6__6__0_ccff_tail));

	sb_10__0_ sb_10__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__20_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__18_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_16_ccff_tail),
		.chany_top_out(sb_10__0__0_chany_top_out[0:104]),
		.chanx_left_out(sb_10__0__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__0__0_ccff_tail));

	sb_10__1_ sb_10__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__21_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__20_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_9_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__19_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_18_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_18_ccff_tail),
		.chany_top_out(sb_10__1__0_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__1__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__1__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__1__0_ccff_tail));

	sb_10__2_ sb_10__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_0__1__21_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_8_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__2__9_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_71_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_19_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_63_ccff_tail),
		.chany_top_out(sb_10__2__0_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__2__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__2__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__2__0_ccff_tail));

	sb_10__3_ sb_10__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__1_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_7_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_71_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__61_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_72_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_71_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_71_ccff_tail),
		.chany_top_out(sb_10__3__0_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__3__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__3__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__3__0_ccff_tail));

	sb_10__3_ sb_10__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__2_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__1_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_6_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_72_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__62_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_73_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_72_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_65_ccff_tail),
		.chany_top_out(sb_10__3__1_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__3__1_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__3__1_chanx_left_out[0:104]),
		.ccff_tail(sb_10__3__1_ccff_tail));

	sb_10__3_ sb_10__7_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__4_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__3_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__63_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_75_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_74_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_74_ccff_tail),
		.chany_top_out(sb_10__3__2_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__3__2_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__3__2_chanx_left_out[0:104]),
		.ccff_tail(sb_10__3__2_ccff_tail));

	sb_10__3_ sb_10__8_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__5_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__4_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_75_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__64_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_76_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_75_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_69_ccff_tail),
		.chany_top_out(sb_10__3__3_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__3__3_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__3__3_chanx_left_out[0:104]),
		.ccff_tail(sb_10__3__3_ccff_tail));

	sb_10__3_ sb_10__9_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__6_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__5_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_76_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__65_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_77_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_76_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_76_ccff_tail),
		.chany_top_out(sb_10__3__4_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__3__4_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__3__4_chanx_left_out[0:104]),
		.ccff_tail(sb_10__3__4_ccff_tail));

	sb_10__5_ sb_10__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__6__0_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__3__2_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_73_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_6__5__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_0_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_5_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_9_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_13_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_17_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_21_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_25_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_29_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_1_33_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_6_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_10_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_14_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_18_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_22_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_26_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_30_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_2_34_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_3_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_7_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_11_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_15_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_19_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_23_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_27_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_3_31_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_odata_4_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_oack_3_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_1_1_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_olck_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_73_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_73_ccff_tail),
		.chany_top_out(sb_10__5__0_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__5__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__5__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__5__0_ccff_tail));

	sb_10__6_ sb_10__6_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_10__3__3_chany_bottom_out[0:104]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_74_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_10__6__0_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_0_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_0_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_4_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_4_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_8_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_12_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_16_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_16_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_20_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_20_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_24_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_24_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_28_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_28_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_1_32_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_1_32_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_1_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_5_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_9_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_13_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_17_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_17_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_21_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_21_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_25_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_25_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_29_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_29_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_2_33_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_2_33_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_2_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_2_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_6_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_6_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_10_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_14_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_18_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_18_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_22_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_22_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_26_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_26_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_30_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_30_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_3_34_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_3_34_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_odata_4_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_odata_4_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovalid_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ovch_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_oack_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_oack_3_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_0_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_0_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_2_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_2_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_ordy_4_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_ordy_4_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_1_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_1_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_olck_3_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_olck_3_0_),
		.chanx_left_in(cbx_6__6__1_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_74_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_0_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_0_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_3_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_7_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_7_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_11_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_11_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_15_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_15_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_19_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_19_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_23_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_23_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_27_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_27_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_1_31_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_1_31_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_4_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_8_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_12_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_12_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_16_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_16_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_20_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_20_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_24_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_24_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_28_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_28_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_2_32_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_2_32_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_5_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_9_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_9_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_13_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_13_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_17_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_17_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_21_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_21_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_25_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_25_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_29_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_29_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_3_33_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_3_33_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_odata_4_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_odata_4_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovalid_3_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ovch_2_0_(grid_router_1_top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_oack_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_oack_4_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_1_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_1_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_ordy_3_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_ordy_3_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_0_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_0_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_2_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_2_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_olck_4_1_(grid_router_1_top_width_0_height_0_subtile_0__pin_olck_4_1_),
		.ccff_head(grid_clb_67_ccff_tail),
		.chany_top_out(sb_10__6__0_chany_top_out[0:104]),
		.chany_bottom_out(sb_10__6__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__6__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__6__0_ccff_tail));

	sb_10__10_ sb_10__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_10__3__6_chany_top_out[0:104]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_77_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__10__9_chanx_right_out[0:104]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_9_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_77_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_10__10__0_chany_bottom_out[0:104]),
		.chanx_left_out(sb_10__10__0_chanx_left_out[0:104]),
		.ccff_tail(sb_10__10__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_1__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_2__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_3__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__6_ccff_tail));

	cbx_1__0_ cbx_4__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__7_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__8_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__8_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__8_ccff_tail));

	cbx_1__0_ cbx_5__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__0__9_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__9_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__9_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__5_ccff_tail),
		.chanx_left_out(cbx_1__0__10_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__10_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__10_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__10_ccff_tail));

	cbx_1__0_ cbx_6__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__0__11_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__11_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__11_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__11_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__6_ccff_tail),
		.chanx_left_out(cbx_1__0__12_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__12_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__12_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__12_ccff_tail));

	cbx_1__0_ cbx_7__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__0__13_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__13_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__13_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__13_ccff_tail));

	cbx_1__0_ cbx_8__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__7_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__7_ccff_tail),
		.chanx_left_out(cbx_1__0__14_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__14_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__14_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__14_ccff_tail));

	cbx_1__0_ cbx_8__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__0__15_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__15_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__15_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__15_ccff_tail));

	cbx_1__0_ cbx_9__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__7_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__0__8_chanx_left_out[0:104]),
		.ccff_head(sb_1__0__8_ccff_tail),
		.chanx_left_out(cbx_1__0__16_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__16_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__16_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__16_ccff_tail));

	cbx_1__0_ cbx_9__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:104]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__0__17_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__17_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__17_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__17_ccff_tail));

	cbx_1__0_ cbx_10__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__8_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__0__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__18_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__18_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__18_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__18_ccff_tail));

	cbx_1__0_ cbx_10__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__1__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__1__0_ccff_tail),
		.chanx_left_out(cbx_1__0__19_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__0__19_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__19_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__19_ccff_tail));

	cbx_1__2_ cbx_1__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__0_ccff_tail));

	cbx_1__2_ cbx_2__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__1_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__1_ccff_tail),
		.chanx_left_out(cbx_1__2__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__1_ccff_tail));

	cbx_1__2_ cbx_3__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__2_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__2_ccff_tail),
		.chanx_left_out(cbx_1__2__2_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__2_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__2_ccff_tail));

	cbx_1__2_ cbx_4__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__3_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__3_ccff_tail),
		.chanx_left_out(cbx_1__2__3_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__3_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__3_ccff_tail));

	cbx_1__2_ cbx_5__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__4_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__4_ccff_tail),
		.chanx_left_out(cbx_1__2__4_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__4_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__4_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__4_ccff_tail));

	cbx_1__2_ cbx_6__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__5_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__5_ccff_tail),
		.chanx_left_out(cbx_1__2__5_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__5_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__5_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__5_ccff_tail));

	cbx_1__2_ cbx_7__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__6_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__6_ccff_tail),
		.chanx_left_out(cbx_1__2__6_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__6_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__6_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__6_ccff_tail));

	cbx_1__2_ cbx_8__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__7_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__7_ccff_tail),
		.chanx_left_out(cbx_1__2__7_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__7_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__7_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__7_ccff_tail));

	cbx_1__2_ cbx_9__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__7_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__2__8_chanx_left_out[0:104]),
		.ccff_head(sb_1__2__8_ccff_tail),
		.chanx_left_out(cbx_1__2__8_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__8_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__8_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__8_ccff_tail));

	cbx_1__2_ cbx_10__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__8_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__2__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__9_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__2__9_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__2__9_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__2__9_ccff_tail));

	cbx_1__3_ cbx_1__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__0_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__0_ccff_tail));

	cbx_1__3_ cbx_1__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__1_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__1_ccff_tail),
		.chanx_left_out(cbx_1__3__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__1_ccff_tail));

	cbx_1__3_ cbx_1__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__2_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__2_ccff_tail),
		.chanx_left_out(cbx_1__3__2_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__2_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__2_ccff_tail));

	cbx_1__3_ cbx_1__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__3_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__3_ccff_tail),
		.chanx_left_out(cbx_1__3__3_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__3_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__3_ccff_tail));

	cbx_1__3_ cbx_1__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__4_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__4_ccff_tail),
		.chanx_left_out(cbx_1__3__4_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__4_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__4_ccff_tail));

	cbx_1__3_ cbx_1__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__5_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__5_ccff_tail),
		.chanx_left_out(cbx_1__3__5_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__5_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__5_ccff_tail));

	cbx_1__3_ cbx_1__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__6_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__6_ccff_tail),
		.chanx_left_out(cbx_1__3__6_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__6_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__6_ccff_tail));

	cbx_1__3_ cbx_2__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__7_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__7_ccff_tail),
		.chanx_left_out(cbx_1__3__7_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__7_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__7_ccff_tail));

	cbx_1__3_ cbx_2__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__8_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__8_ccff_tail),
		.chanx_left_out(cbx_1__3__8_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__8_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__8_ccff_tail));

	cbx_1__3_ cbx_2__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__9_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__9_ccff_tail),
		.chanx_left_out(cbx_1__3__9_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__9_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__9_ccff_tail));

	cbx_1__3_ cbx_2__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__10_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__10_ccff_tail),
		.chanx_left_out(cbx_1__3__10_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__10_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__10_ccff_tail));

	cbx_1__3_ cbx_2__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__11_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__11_ccff_tail),
		.chanx_left_out(cbx_1__3__11_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__11_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__11_ccff_tail));

	cbx_1__3_ cbx_2__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__12_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__12_ccff_tail),
		.chanx_left_out(cbx_1__3__12_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__12_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__12_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__12_ccff_tail));

	cbx_1__3_ cbx_2__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__13_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__13_ccff_tail),
		.chanx_left_out(cbx_1__3__13_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__13_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__13_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__13_ccff_tail));

	cbx_1__3_ cbx_3__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__7_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__14_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__14_ccff_tail),
		.chanx_left_out(cbx_1__3__14_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__14_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__14_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__14_ccff_tail));

	cbx_1__3_ cbx_3__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__8_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__15_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__15_ccff_tail),
		.chanx_left_out(cbx_1__3__15_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__15_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__15_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__15_ccff_tail));

	cbx_1__3_ cbx_3__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__9_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__16_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__16_ccff_tail),
		.chanx_left_out(cbx_1__3__16_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__16_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__16_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__16_ccff_tail));

	cbx_1__3_ cbx_3__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__10_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__17_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__17_ccff_tail),
		.chanx_left_out(cbx_1__3__17_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__17_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__17_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__17_ccff_tail));

	cbx_1__3_ cbx_3__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__11_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__18_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__18_ccff_tail),
		.chanx_left_out(cbx_1__3__18_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__18_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__18_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__18_ccff_tail));

	cbx_1__3_ cbx_3__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__12_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__19_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__19_ccff_tail),
		.chanx_left_out(cbx_1__3__19_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__19_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__19_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__19_ccff_tail));

	cbx_1__3_ cbx_3__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__13_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__20_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__20_ccff_tail),
		.chanx_left_out(cbx_1__3__20_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__20_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__20_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__20_ccff_tail));

	cbx_1__3_ cbx_4__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__14_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__21_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__21_ccff_tail),
		.chanx_left_out(cbx_1__3__21_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__21_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__21_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__21_ccff_tail));

	cbx_1__3_ cbx_4__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__15_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__22_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__22_ccff_tail),
		.chanx_left_out(cbx_1__3__22_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__22_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__22_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__22_ccff_tail));

	cbx_1__3_ cbx_4__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__16_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__23_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__23_ccff_tail),
		.chanx_left_out(cbx_1__3__23_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__23_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__23_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__23_ccff_tail));

	cbx_1__3_ cbx_4__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__17_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__24_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__24_ccff_tail),
		.chanx_left_out(cbx_1__3__24_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__24_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__24_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__24_ccff_tail));

	cbx_1__3_ cbx_4__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__18_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__25_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__25_ccff_tail),
		.chanx_left_out(cbx_1__3__25_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__25_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__25_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__25_ccff_tail));

	cbx_1__3_ cbx_4__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__19_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__26_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__26_ccff_tail),
		.chanx_left_out(cbx_1__3__26_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__26_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__26_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__26_ccff_tail));

	cbx_1__3_ cbx_4__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__20_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__27_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__27_ccff_tail),
		.chanx_left_out(cbx_1__3__27_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__27_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__27_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__27_ccff_tail));

	cbx_1__3_ cbx_5__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__21_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__28_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__28_ccff_tail),
		.chanx_left_out(cbx_1__3__28_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__28_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__28_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__28_ccff_tail));

	cbx_1__3_ cbx_5__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__22_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__29_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__29_ccff_tail),
		.chanx_left_out(cbx_1__3__29_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__29_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__29_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__29_ccff_tail));

	cbx_1__3_ cbx_5__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__23_chanx_right_out[0:104]),
		.chanx_right_in(sb_5__5__0_chanx_left_out[0:104]),
		.ccff_head(sb_5__5__0_ccff_tail),
		.chanx_left_out(cbx_1__3__30_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__30_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__30_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__30_ccff_tail));

	cbx_1__3_ cbx_5__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__24_chanx_right_out[0:104]),
		.chanx_right_in(sb_5__6__0_chanx_left_out[0:104]),
		.ccff_head(sb_5__6__0_ccff_tail),
		.chanx_left_out(cbx_1__3__31_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__31_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__31_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__31_ccff_tail));

	cbx_1__3_ cbx_5__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__25_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__30_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__30_ccff_tail),
		.chanx_left_out(cbx_1__3__32_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__32_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__32_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__32_ccff_tail));

	cbx_1__3_ cbx_5__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__26_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__31_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__31_ccff_tail),
		.chanx_left_out(cbx_1__3__33_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__33_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__33_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__33_ccff_tail));

	cbx_1__3_ cbx_5__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__27_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__32_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__32_ccff_tail),
		.chanx_left_out(cbx_1__3__34_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__34_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__34_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__34_ccff_tail));

	cbx_1__3_ cbx_6__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__28_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__33_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__33_ccff_tail),
		.chanx_left_out(cbx_1__3__35_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__35_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__35_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__35_ccff_tail));

	cbx_1__3_ cbx_6__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__29_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__34_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__34_ccff_tail),
		.chanx_left_out(cbx_1__3__36_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__36_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__36_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__36_ccff_tail));

	cbx_1__3_ cbx_6__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__30_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__35_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__35_ccff_tail),
		.chanx_left_out(cbx_1__3__37_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__37_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__37_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__37_ccff_tail));

	cbx_1__3_ cbx_6__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__31_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__36_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__36_ccff_tail),
		.chanx_left_out(cbx_1__3__38_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__38_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__38_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__38_ccff_tail));

	cbx_1__3_ cbx_6__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__32_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__37_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__37_ccff_tail),
		.chanx_left_out(cbx_1__3__39_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__39_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__39_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__39_ccff_tail));

	cbx_1__3_ cbx_7__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__33_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__38_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__38_ccff_tail),
		.chanx_left_out(cbx_1__3__40_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__40_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__40_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__40_ccff_tail));

	cbx_1__3_ cbx_7__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__34_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__39_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__39_ccff_tail),
		.chanx_left_out(cbx_1__3__41_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__41_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__41_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__41_ccff_tail));

	cbx_1__3_ cbx_7__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_6__5__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__40_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__40_ccff_tail),
		.chanx_left_out(cbx_1__3__42_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__42_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__42_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__42_ccff_tail));

	cbx_1__3_ cbx_7__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_6__6__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__41_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__41_ccff_tail),
		.chanx_left_out(cbx_1__3__43_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__43_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__43_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__43_ccff_tail));

	cbx_1__3_ cbx_7__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__35_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__42_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__42_ccff_tail),
		.chanx_left_out(cbx_1__3__44_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__44_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__44_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__44_ccff_tail));

	cbx_1__3_ cbx_7__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__36_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__43_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__43_ccff_tail),
		.chanx_left_out(cbx_1__3__45_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__45_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__45_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__45_ccff_tail));

	cbx_1__3_ cbx_7__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__37_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__44_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__44_ccff_tail),
		.chanx_left_out(cbx_1__3__46_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__46_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__46_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__46_ccff_tail));

	cbx_1__3_ cbx_8__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__38_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__45_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__45_ccff_tail),
		.chanx_left_out(cbx_1__3__47_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__47_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__47_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__47_ccff_tail));

	cbx_1__3_ cbx_8__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__39_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__46_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__46_ccff_tail),
		.chanx_left_out(cbx_1__3__48_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__48_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__48_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__48_ccff_tail));

	cbx_1__3_ cbx_8__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__40_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__47_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__47_ccff_tail),
		.chanx_left_out(cbx_1__3__49_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__49_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__49_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__49_ccff_tail));

	cbx_1__3_ cbx_8__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__41_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__48_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__48_ccff_tail),
		.chanx_left_out(cbx_1__3__50_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__50_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__50_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__50_ccff_tail));

	cbx_1__3_ cbx_8__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__42_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__49_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__49_ccff_tail),
		.chanx_left_out(cbx_1__3__51_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__51_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__51_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__51_ccff_tail));

	cbx_1__3_ cbx_8__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__43_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__50_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__50_ccff_tail),
		.chanx_left_out(cbx_1__3__52_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__52_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__52_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__52_ccff_tail));

	cbx_1__3_ cbx_8__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__44_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__51_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__51_ccff_tail),
		.chanx_left_out(cbx_1__3__53_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__53_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__53_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__53_ccff_tail));

	cbx_1__3_ cbx_9__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__45_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__52_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__52_ccff_tail),
		.chanx_left_out(cbx_1__3__54_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__54_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__54_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__54_ccff_tail));

	cbx_1__3_ cbx_9__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__46_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__53_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__53_ccff_tail),
		.chanx_left_out(cbx_1__3__55_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__55_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__55_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__55_ccff_tail));

	cbx_1__3_ cbx_9__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__47_chanx_right_out[0:104]),
		.chanx_right_in(sb_5__5__1_chanx_left_out[0:104]),
		.ccff_head(sb_5__5__1_ccff_tail),
		.chanx_left_out(cbx_1__3__56_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__56_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__56_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__56_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__56_ccff_tail));

	cbx_1__3_ cbx_9__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__48_chanx_right_out[0:104]),
		.chanx_right_in(sb_5__6__1_chanx_left_out[0:104]),
		.ccff_head(sb_5__6__1_ccff_tail),
		.chanx_left_out(cbx_1__3__57_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__57_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__57_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__57_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__57_ccff_tail));

	cbx_1__3_ cbx_9__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__49_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__54_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__54_ccff_tail),
		.chanx_left_out(cbx_1__3__58_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__58_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__58_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__58_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__58_ccff_tail));

	cbx_1__3_ cbx_9__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__50_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__55_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__55_ccff_tail),
		.chanx_left_out(cbx_1__3__59_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__59_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__59_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__59_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__59_ccff_tail));

	cbx_1__3_ cbx_9__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__51_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__3__56_chanx_left_out[0:104]),
		.ccff_head(sb_1__3__56_ccff_tail),
		.chanx_left_out(cbx_1__3__60_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__60_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__60_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__60_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__60_ccff_tail));

	cbx_1__3_ cbx_10__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__52_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__3__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__61_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__61_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__61_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__61_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__61_ccff_tail));

	cbx_1__3_ cbx_10__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__53_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__3__1_chanx_left_out[0:104]),
		.ccff_head(sb_10__3__1_ccff_tail),
		.chanx_left_out(cbx_1__3__62_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__62_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__62_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__62_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__62_ccff_tail));

	cbx_1__3_ cbx_10__7_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__54_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__3__2_chanx_left_out[0:104]),
		.ccff_head(sb_10__3__2_ccff_tail),
		.chanx_left_out(cbx_1__3__63_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__63_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__63_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__63_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__63_ccff_tail));

	cbx_1__3_ cbx_10__8_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__55_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__3__3_chanx_left_out[0:104]),
		.ccff_head(sb_10__3__3_ccff_tail),
		.chanx_left_out(cbx_1__3__64_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__64_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__64_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__64_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__64_ccff_tail));

	cbx_1__3_ cbx_10__9_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__56_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__3__4_chanx_left_out[0:104]),
		.ccff_head(sb_10__3__4_ccff_tail),
		.chanx_left_out(cbx_1__3__65_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__3__65_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__65_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__65_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__65_ccff_tail));

	cbx_1__10_ cbx_1__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__10__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__0_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__0_ccff_tail),
		.chanx_left_out(cbx_1__10__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__0_ccff_tail));

	cbx_1__10_ cbx_2__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__1_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__1_ccff_tail),
		.chanx_left_out(cbx_1__10__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__1_ccff_tail));

	cbx_1__10_ cbx_3__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__2_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__2_ccff_tail),
		.chanx_left_out(cbx_1__10__2_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__2_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__2_ccff_tail));

	cbx_1__10_ cbx_4__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__2_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__3_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__3_ccff_tail),
		.chanx_left_out(cbx_1__10__3_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__3_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__3_ccff_tail));

	cbx_1__10_ cbx_5__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__3_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__4_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__4_ccff_tail),
		.chanx_left_out(cbx_1__10__4_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__4_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__4_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__4_ccff_tail));

	cbx_1__10_ cbx_6__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__4_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__5_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__5_ccff_tail),
		.chanx_left_out(cbx_1__10__5_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__5_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__5_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__5_ccff_tail));

	cbx_1__10_ cbx_7__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__5_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__6_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__6_ccff_tail),
		.chanx_left_out(cbx_1__10__6_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__6_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__6_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__6_ccff_tail));

	cbx_1__10_ cbx_8__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__6_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__7_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__7_ccff_tail),
		.chanx_left_out(cbx_1__10__7_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__7_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__7_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__7_ccff_tail));

	cbx_1__10_ cbx_9__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__7_chanx_right_out[0:104]),
		.chanx_right_in(sb_1__10__8_chanx_left_out[0:104]),
		.ccff_head(sb_1__10__8_ccff_tail),
		.chanx_left_out(cbx_1__10__8_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__8_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__8_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__8_ccff_tail));

	cbx_1__10_ cbx_10__10_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__10__8_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__10__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__10__0_ccff_tail),
		.chanx_left_out(cbx_1__10__9_chanx_left_out[0:104]),
		.chanx_right_out(cbx_1__10__9_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__10__9_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__10__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__10__9_ccff_tail));

	cbx_6__5_ cbx_6__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_5__5__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_6__5__0_chanx_left_out[0:104]),
		.ccff_head(sb_6__5__0_ccff_tail),
		.chanx_left_out(cbx_6__5__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_6__5__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_6__5__0_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_6__5__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_6__5__0_ccff_tail));

	cbx_6__5_ cbx_10__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_5__5__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__5__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__5__0_ccff_tail),
		.chanx_left_out(cbx_6__5__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_6__5__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_my_xpos_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_0_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_1_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_2_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_4_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_8_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_12_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_16_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_20_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_24_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_28_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_3_32_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_9_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_13_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_17_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_21_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_25_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_29_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_idata_4_33_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_0_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_2_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_iack_4_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_1_0_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_(cbx_6__5__1_top_grid_bottom_width_0_height_0_subtile_0__pin_ilck_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_6__5__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_6__5__1_ccff_tail));

	cbx_6__6_ cbx_6__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_5__6__0_chanx_right_out[0:104]),
		.chanx_right_in(sb_6__6__0_chanx_left_out[0:104]),
		.ccff_head(sb_6__6__0_ccff_tail),
		.chanx_left_out(cbx_6__6__0_chanx_left_out[0:104]),
		.chanx_right_out(cbx_6__6__0_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_6__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_6__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_6__6__0_ccff_tail));

	cbx_6__6_ cbx_10__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_5__6__1_chanx_right_out[0:104]),
		.chanx_right_in(sb_10__6__0_chanx_left_out[0:104]),
		.ccff_head(sb_10__6__0_ccff_tail),
		.chanx_left_out(cbx_6__6__1_chanx_left_out[0:104]),
		.chanx_right_out(cbx_6__6__1_chanx_right_out[0:104]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_6__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_rst__0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_my_ypos_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_0_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_1_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_2_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_2_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_10_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_14_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_18_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_22_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_26_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_30_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_3_34_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_11_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_15_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_19_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_23_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_27_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_idata_4_31_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_iack_3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_(cbx_6__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_ilck_4_0_),
		.ccff_tail(cbx_6__6__1_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:104]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:104]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:104]),
		.chany_top_in(sb_0__2__0_chany_bottom_out[0:104]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_1__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_1__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_2__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__1_ cby_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__5_ccff_tail));

	cby_0__1_ cby_3__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__6_ccff_tail));

	cby_0__1_ cby_3__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__2_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__7_ccff_tail));

	cby_0__1_ cby_4__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__6_ccff_tail),
		.chany_bottom_out(cby_0__1__8_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__8_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__8_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__8_ccff_tail));

	cby_0__1_ cby_4__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__3_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__7_ccff_tail),
		.chany_bottom_out(cby_0__1__9_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__9_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__9_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__9_ccff_tail));

	cby_0__1_ cby_5__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__8_ccff_tail),
		.chany_bottom_out(cby_0__1__10_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__10_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__10_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__10_ccff_tail));

	cby_0__1_ cby_5__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__4_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__9_ccff_tail),
		.chany_bottom_out(cby_0__1__11_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__11_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__11_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__11_ccff_tail));

	cby_0__1_ cby_6__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__10_ccff_tail),
		.chany_bottom_out(cby_0__1__12_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__12_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__12_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__12_ccff_tail));

	cby_0__1_ cby_6__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__5_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__11_ccff_tail),
		.chany_bottom_out(cby_0__1__13_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__13_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__13_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__13_ccff_tail));

	cby_0__1_ cby_7__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__12_ccff_tail),
		.chany_bottom_out(cby_0__1__14_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__14_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__14_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__14_ccff_tail));

	cby_0__1_ cby_7__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__6_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__13_ccff_tail),
		.chany_bottom_out(cby_0__1__15_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__15_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__15_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__15_ccff_tail));

	cby_0__1_ cby_8__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__7_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__14_ccff_tail),
		.chany_bottom_out(cby_0__1__16_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__16_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__16_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__16_ccff_tail));

	cby_0__1_ cby_8__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__7_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__15_ccff_tail),
		.chany_bottom_out(cby_0__1__17_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__17_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__17_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__17_ccff_tail));

	cby_0__1_ cby_9__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__8_chany_top_out[0:104]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__16_ccff_tail),
		.chany_bottom_out(cby_0__1__18_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__18_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__18_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__18_ccff_tail));

	cby_0__1_ cby_9__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:104]),
		.chany_top_in(sb_1__2__8_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__17_ccff_tail),
		.chany_bottom_out(cby_0__1__19_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__19_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__19_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__19_ccff_tail));

	cby_0__1_ cby_10__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__0__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__1__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__18_ccff_tail),
		.chany_bottom_out(cby_0__1__20_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__20_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__20_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__20_ccff_tail));

	cby_0__1_ cby_10__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__1__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__2__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__0__19_ccff_tail),
		.chany_bottom_out(cby_0__1__21_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__1__21_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__21_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__21_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__21_ccff_tail));

	cby_0__3_ cby_0__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__2__0_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__0_chany_bottom_out[0:104]),
		.ccff_head(sb_0__2__0_ccff_tail),
		.chany_bottom_out(cby_0__3__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__0_ccff_tail));

	cby_0__3_ cby_0__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__0_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__1_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__0_ccff_tail),
		.chany_bottom_out(cby_0__3__1_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__1_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__1_ccff_tail));

	cby_0__3_ cby_0__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__1_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__2_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__1_ccff_tail),
		.chany_bottom_out(cby_0__3__2_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__2_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__2_ccff_tail));

	cby_0__3_ cby_0__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__2_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__3_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__2_ccff_tail),
		.chany_bottom_out(cby_0__3__3_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__3_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__3_ccff_tail));

	cby_0__3_ cby_0__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__3_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__4_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__3_ccff_tail),
		.chany_bottom_out(cby_0__3__4_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__4_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__4_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__4_ccff_tail));

	cby_0__3_ cby_0__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__4_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__5_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__4_ccff_tail),
		.chany_bottom_out(cby_0__3__5_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__5_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__5_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__5_ccff_tail));

	cby_0__3_ cby_0__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__5_chany_top_out[0:104]),
		.chany_top_in(sb_0__3__6_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__5_ccff_tail),
		.chany_bottom_out(cby_0__3__6_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__6_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__6_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__6_ccff_tail));

	cby_0__3_ cby_0__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__6_chany_top_out[0:104]),
		.chany_top_in(sb_0__10__0_chany_bottom_out[0:104]),
		.ccff_head(sb_0__3__6_ccff_tail),
		.chany_bottom_out(cby_0__3__7_chany_bottom_out[0:104]),
		.chany_top_out(cby_0__3__7_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__3__7_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__3__7_ccff_tail));

	cby_1__3_ cby_1__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__0_ccff_tail),
		.chany_bottom_out(cby_1__3__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__0_ccff_tail));

	cby_1__3_ cby_1__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__0_ccff_tail),
		.chany_bottom_out(cby_1__3__1_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__1_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__1_ccff_tail));

	cby_1__3_ cby_1__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__1_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__2_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__1_ccff_tail),
		.chany_bottom_out(cby_1__3__2_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__2_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__2_ccff_tail));

	cby_1__3_ cby_1__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__2_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__3_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__2_ccff_tail),
		.chany_bottom_out(cby_1__3__3_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__3_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__3_ccff_tail));

	cby_1__3_ cby_1__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__3_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__4_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__3_ccff_tail),
		.chany_bottom_out(cby_1__3__4_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__4_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__4_ccff_tail));

	cby_1__3_ cby_1__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__4_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__5_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__4_ccff_tail),
		.chany_bottom_out(cby_1__3__5_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__5_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__5_ccff_tail));

	cby_1__3_ cby_1__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__5_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__6_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__5_ccff_tail),
		.chany_bottom_out(cby_1__3__6_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__6_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__6_ccff_tail));

	cby_1__3_ cby_1__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__6_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__6_ccff_tail),
		.chany_bottom_out(cby_1__3__7_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__7_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__7_ccff_tail));

	cby_1__3_ cby_2__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__1_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__7_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__1_ccff_tail),
		.chany_bottom_out(cby_1__3__8_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__8_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__8_ccff_tail));

	cby_1__3_ cby_2__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__7_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__8_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__7_ccff_tail),
		.chany_bottom_out(cby_1__3__9_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__9_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__9_ccff_tail));

	cby_1__3_ cby_2__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__8_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__9_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__8_ccff_tail),
		.chany_bottom_out(cby_1__3__10_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__10_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__10_ccff_tail));

	cby_1__3_ cby_2__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__9_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__10_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__9_ccff_tail),
		.chany_bottom_out(cby_1__3__11_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__11_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__11_ccff_tail));

	cby_1__3_ cby_2__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__10_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__11_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__10_ccff_tail),
		.chany_bottom_out(cby_1__3__12_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__12_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__12_ccff_tail));

	cby_1__3_ cby_2__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__11_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__12_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__11_ccff_tail),
		.chany_bottom_out(cby_1__3__13_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__13_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__13_ccff_tail));

	cby_1__3_ cby_2__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__12_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__13_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__12_ccff_tail),
		.chany_bottom_out(cby_1__3__14_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__14_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__14_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__14_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__14_ccff_tail));

	cby_1__3_ cby_2__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__13_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__13_ccff_tail),
		.chany_bottom_out(cby_1__3__15_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__15_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__15_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__15_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__15_ccff_tail));

	cby_1__3_ cby_3__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__2_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__14_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__2_ccff_tail),
		.chany_bottom_out(cby_1__3__16_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__16_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__16_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__16_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__16_ccff_tail));

	cby_1__3_ cby_3__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__14_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__15_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__14_ccff_tail),
		.chany_bottom_out(cby_1__3__17_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__17_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__17_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__17_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__17_ccff_tail));

	cby_1__3_ cby_3__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__15_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__16_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__15_ccff_tail),
		.chany_bottom_out(cby_1__3__18_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__18_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__18_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__18_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__18_ccff_tail));

	cby_1__3_ cby_3__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__16_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__17_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__16_ccff_tail),
		.chany_bottom_out(cby_1__3__19_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__19_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__19_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__19_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__19_ccff_tail));

	cby_1__3_ cby_3__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__17_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__18_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__17_ccff_tail),
		.chany_bottom_out(cby_1__3__20_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__20_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__20_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__20_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__20_ccff_tail));

	cby_1__3_ cby_3__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__18_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__19_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__18_ccff_tail),
		.chany_bottom_out(cby_1__3__21_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__21_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__21_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__21_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__21_ccff_tail));

	cby_1__3_ cby_3__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__19_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__20_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__19_ccff_tail),
		.chany_bottom_out(cby_1__3__22_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__22_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__22_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__22_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__22_ccff_tail));

	cby_1__3_ cby_3__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__20_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__2_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__20_ccff_tail),
		.chany_bottom_out(cby_1__3__23_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__23_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__23_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__23_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__23_ccff_tail));

	cby_1__3_ cby_4__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__3_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__21_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__3_ccff_tail),
		.chany_bottom_out(cby_1__3__24_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__24_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__24_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__24_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__24_ccff_tail));

	cby_1__3_ cby_4__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__21_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__22_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__21_ccff_tail),
		.chany_bottom_out(cby_1__3__25_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__25_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__25_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__25_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__25_ccff_tail));

	cby_1__3_ cby_4__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__22_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__23_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__22_ccff_tail),
		.chany_bottom_out(cby_1__3__26_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__26_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__26_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__26_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__26_ccff_tail));

	cby_1__3_ cby_4__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__23_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__24_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__23_ccff_tail),
		.chany_bottom_out(cby_1__3__27_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__27_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__27_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__27_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__27_ccff_tail));

	cby_1__3_ cby_4__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__24_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__25_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__24_ccff_tail),
		.chany_bottom_out(cby_1__3__28_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__28_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__28_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__28_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__28_ccff_tail));

	cby_1__3_ cby_4__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__25_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__26_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__25_ccff_tail),
		.chany_bottom_out(cby_1__3__29_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__29_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__29_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__29_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__29_ccff_tail));

	cby_1__3_ cby_4__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__26_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__27_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__26_ccff_tail),
		.chany_bottom_out(cby_1__3__30_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__30_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__30_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__30_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__30_ccff_tail));

	cby_1__3_ cby_4__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__27_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__3_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__27_ccff_tail),
		.chany_bottom_out(cby_1__3__31_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__31_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__31_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__31_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__31_ccff_tail));

	cby_1__3_ cby_5__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__4_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__28_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__4_ccff_tail),
		.chany_bottom_out(cby_1__3__32_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__32_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__32_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__32_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__32_ccff_tail));

	cby_1__3_ cby_5__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__28_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__29_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__28_ccff_tail),
		.chany_bottom_out(cby_1__3__33_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__33_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__33_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__33_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__33_ccff_tail));

	cby_1__3_ cby_5__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__29_chany_top_out[0:104]),
		.chany_top_in(sb_5__5__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__29_ccff_tail),
		.chany_bottom_out(cby_1__3__34_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__34_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__34_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__34_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__34_ccff_tail));

	cby_1__3_ cby_5__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__6__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__30_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__31_ccff_tail),
		.chany_bottom_out(cby_1__3__35_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__35_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__35_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__35_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__35_ccff_tail));

	cby_1__3_ cby_5__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__30_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__31_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__32_ccff_tail),
		.chany_bottom_out(cby_1__3__36_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__36_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__36_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__36_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__36_ccff_tail));

	cby_1__3_ cby_5__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__31_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__32_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__33_ccff_tail),
		.chany_bottom_out(cby_1__3__37_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__37_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__37_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__37_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__37_ccff_tail));

	cby_1__3_ cby_5__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__32_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__4_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__34_ccff_tail),
		.chany_bottom_out(cby_1__3__38_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__38_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__38_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__38_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__38_ccff_tail));

	cby_1__3_ cby_6__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__5_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__33_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__5_ccff_tail),
		.chany_bottom_out(cby_1__3__39_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__39_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__39_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__39_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__39_ccff_tail));

	cby_1__3_ cby_6__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__33_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__34_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__35_ccff_tail),
		.chany_bottom_out(cby_1__3__40_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__40_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__40_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__40_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__40_ccff_tail));

	cby_1__3_ cby_6__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__34_chany_top_out[0:104]),
		.chany_top_in(sb_6__5__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__36_ccff_tail),
		.chany_bottom_out(cby_1__3__41_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__41_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__41_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__41_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__41_ccff_tail));

	cby_1__3_ cby_6__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__6__0_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__35_chany_bottom_out[0:104]),
		.ccff_head(cbx_6__6__0_ccff_tail),
		.chany_bottom_out(cby_1__3__42_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__42_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__42_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__42_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__42_ccff_tail));

	cby_1__3_ cby_6__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__35_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__36_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__37_ccff_tail),
		.chany_bottom_out(cby_1__3__43_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__43_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__43_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__43_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__43_ccff_tail));

	cby_1__3_ cby_6__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__36_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__37_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__38_ccff_tail),
		.chany_bottom_out(cby_1__3__44_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__44_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__44_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__44_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__44_ccff_tail));

	cby_1__3_ cby_6__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__37_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__5_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__39_ccff_tail),
		.chany_bottom_out(cby_1__3__45_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__45_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__45_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__45_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__45_ccff_tail));

	cby_1__3_ cby_7__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__6_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__38_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__6_ccff_tail),
		.chany_bottom_out(cby_1__3__46_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__46_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__46_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__46_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__46_ccff_tail));

	cby_1__3_ cby_7__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__38_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__39_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__40_ccff_tail),
		.chany_bottom_out(cby_1__3__47_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__47_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__47_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__47_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__47_ccff_tail));

	cby_1__3_ cby_7__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__39_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__40_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__41_ccff_tail),
		.chany_bottom_out(cby_1__3__48_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__48_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__48_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__48_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__48_ccff_tail));

	cby_1__3_ cby_7__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__40_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__41_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__42_ccff_tail),
		.chany_bottom_out(cby_1__3__49_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__49_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__49_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__49_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__49_ccff_tail));

	cby_1__3_ cby_7__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__41_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__42_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__43_ccff_tail),
		.chany_bottom_out(cby_1__3__50_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__50_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__50_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__50_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__50_ccff_tail));

	cby_1__3_ cby_7__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__42_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__43_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__44_ccff_tail),
		.chany_bottom_out(cby_1__3__51_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__51_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__51_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__51_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__51_ccff_tail));

	cby_1__3_ cby_7__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__43_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__44_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__45_ccff_tail),
		.chany_bottom_out(cby_1__3__52_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__52_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__52_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__52_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__52_ccff_tail));

	cby_1__3_ cby_7__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__44_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__6_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__46_ccff_tail),
		.chany_bottom_out(cby_1__3__53_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__53_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__53_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__53_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__53_ccff_tail));

	cby_1__3_ cby_8__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__7_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__45_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__7_ccff_tail),
		.chany_bottom_out(cby_1__3__54_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__54_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__54_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__54_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__54_ccff_tail));

	cby_1__3_ cby_8__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__45_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__46_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__47_ccff_tail),
		.chany_bottom_out(cby_1__3__55_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__55_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__55_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__55_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__55_ccff_tail));

	cby_1__3_ cby_8__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__46_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__47_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__48_ccff_tail),
		.chany_bottom_out(cby_1__3__56_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__56_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__56_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__56_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__56_ccff_tail));

	cby_1__3_ cby_8__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__47_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__48_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__49_ccff_tail),
		.chany_bottom_out(cby_1__3__57_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__57_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__57_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__57_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__57_ccff_tail));

	cby_1__3_ cby_8__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__48_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__49_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__50_ccff_tail),
		.chany_bottom_out(cby_1__3__58_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__58_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__58_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__58_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__58_ccff_tail));

	cby_1__3_ cby_8__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__49_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__50_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__51_ccff_tail),
		.chany_bottom_out(cby_1__3__59_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__59_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__59_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__59_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__59_ccff_tail));

	cby_1__3_ cby_8__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__50_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__51_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__52_ccff_tail),
		.chany_bottom_out(cby_1__3__60_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__60_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__60_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__60_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__60_ccff_tail));

	cby_1__3_ cby_8__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__51_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__7_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__53_ccff_tail),
		.chany_bottom_out(cby_1__3__61_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__61_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__61_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__61_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__61_ccff_tail));

	cby_1__3_ cby_9__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__8_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__52_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__8_ccff_tail),
		.chany_bottom_out(cby_1__3__62_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__62_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__62_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__62_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__62_ccff_tail));

	cby_1__3_ cby_9__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__52_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__53_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__54_ccff_tail),
		.chany_bottom_out(cby_1__3__63_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__63_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__63_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__63_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__63_ccff_tail));

	cby_1__3_ cby_9__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__53_chany_top_out[0:104]),
		.chany_top_in(sb_5__5__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__55_ccff_tail),
		.chany_bottom_out(cby_1__3__64_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__64_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__64_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__64_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__64_ccff_tail));

	cby_1__3_ cby_9__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__6__1_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__54_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__57_ccff_tail),
		.chany_bottom_out(cby_1__3__65_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__65_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__65_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__65_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__65_ccff_tail));

	cby_1__3_ cby_9__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__54_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__55_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__58_ccff_tail),
		.chany_bottom_out(cby_1__3__66_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__66_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__66_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__66_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__66_ccff_tail));

	cby_1__3_ cby_9__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__55_chany_top_out[0:104]),
		.chany_top_in(sb_1__3__56_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__59_ccff_tail),
		.chany_bottom_out(cby_1__3__67_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__67_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__67_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__67_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__67_ccff_tail));

	cby_1__3_ cby_9__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__56_chany_top_out[0:104]),
		.chany_top_in(sb_1__10__8_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__60_ccff_tail),
		.chany_bottom_out(cby_1__3__68_chany_bottom_out[0:104]),
		.chany_top_out(cby_1__3__68_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__3__68_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__3__68_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__3__68_ccff_tail));

	cby_5__6_ cby_5__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__5__0_chany_top_out[0:104]),
		.chany_top_in(sb_5__6__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__30_ccff_tail),
		.chany_bottom_out(cby_5__6__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_5__6__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_5__6__0_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__6__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_5__6__0_ccff_tail));

	cby_5__6_ cby_9__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_5__5__1_chany_top_out[0:104]),
		.chany_top_in(sb_5__6__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__56_ccff_tail),
		.chany_bottom_out(cby_5__6__1_chany_bottom_out[0:104]),
		.chany_top_out(cby_5__6__1_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_my_ypos_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_0_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_1_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_2_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_5_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_9_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_13_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_17_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_21_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_25_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_29_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_3_33_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_6_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_10_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_14_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_18_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_22_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_26_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_30_),
		.right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_idata_4_34_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_0_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_2_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_iack_4_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_1_1_),
		.right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_(cby_5__6__1_right_grid_left_width_0_height_0_subtile_0__pin_ilck_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_5__6__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_5__6__1_ccff_tail));

	cby_6__6_ cby_6__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_6__5__0_chany_top_out[0:104]),
		.chany_top_in(sb_6__6__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_6__5__0_ccff_tail),
		.chany_bottom_out(cby_6__6__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_6__6__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_6__6__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_6__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_6__6__0_ccff_tail));

	cby_10__3_ cby_10__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__2__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__3__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__2__9_ccff_tail),
		.chany_bottom_out(cby_10__3__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__0_ccff_tail));

	cby_10__3_ cby_10__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__3__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__3__1_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__61_ccff_tail),
		.chany_bottom_out(cby_10__3__1_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__1_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__1_ccff_tail));

	cby_10__3_ cby_10__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__3__1_chany_top_out[0:104]),
		.chany_top_in(sb_10__5__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__62_ccff_tail),
		.chany_bottom_out(cby_10__3__2_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__2_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__2_ccff_tail));

	cby_10__3_ cby_10__7_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__6__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__3__2_chany_bottom_out[0:104]),
		.ccff_head(cbx_6__6__1_ccff_tail),
		.chany_bottom_out(cby_10__3__3_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__3_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__3_ccff_tail));

	cby_10__3_ cby_10__8_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__3__2_chany_top_out[0:104]),
		.chany_top_in(sb_10__3__3_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__63_ccff_tail),
		.chany_bottom_out(cby_10__3__4_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__4_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__4_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__4_ccff_tail));

	cby_10__3_ cby_10__9_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__3__3_chany_top_out[0:104]),
		.chany_top_in(sb_10__3__4_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__64_ccff_tail),
		.chany_bottom_out(cby_10__3__5_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__5_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__5_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__5_ccff_tail));

	cby_10__3_ cby_10__10_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__3__4_chany_top_out[0:104]),
		.chany_top_in(sb_10__10__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_1__3__65_ccff_tail),
		.chany_bottom_out(cby_10__3__6_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__3__6_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__3__6_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_10__3__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_10__3__6_ccff_tail));

	cby_10__6_ cby_10__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_10__5__0_chany_top_out[0:104]),
		.chany_top_in(sb_10__6__0_chany_bottom_out[0:104]),
		.ccff_head(cbx_6__5__1_ccff_tail),
		.chany_bottom_out(cby_10__6__0_chany_bottom_out[0:104]),
		.chany_top_out(cby_10__6__0_chany_top_out[0:104]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_10__6__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_my_xpos_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_0_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_1_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_2_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_3_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_11_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_15_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_19_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_23_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_27_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_3_31_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_12_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_16_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_20_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_24_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_28_),
		.left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_idata_4_32_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_1_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_iack_3_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_0_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_2_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_(cby_10__6__0_left_grid_right_width_0_height_0_subtile_0__pin_ilck_4_1_),
		.ccff_tail(cby_10__6__0_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




