//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Connection Blocks[1][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Jun 27 10:27:38 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for cby_1__2_ -----
module cby_1__2_(prog_clk,
                 chany_bottom_in,
                 chany_top_in,
                 ccff_head,
                 chany_bottom_out,
                 chany_top_out,
                 right_grid_left_width_0_height_0_subtile_0__pin_I_3_,
                 right_grid_left_width_0_height_0_subtile_0__pin_I_7_,
                 left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_,
                 left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_,
                 left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_,
                 left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_,
                 left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_,
                 ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:188] chany_bottom_in;
//----- INPUT PORTS -----
input [0:188] chany_top_in;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:188] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:188] chany_top_out;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
//----- OUTPUT PORTS -----
output [0:0] right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
//----- OUTPUT PORTS -----
output [0:0] left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:6] mux_tree_tapbuf_size64_0_sram;
wire [0:6] mux_tree_tapbuf_size64_0_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_10_sram;
wire [0:6] mux_tree_tapbuf_size64_10_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_11_sram;
wire [0:6] mux_tree_tapbuf_size64_11_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_12_sram;
wire [0:6] mux_tree_tapbuf_size64_12_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_13_sram;
wire [0:6] mux_tree_tapbuf_size64_13_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_14_sram;
wire [0:6] mux_tree_tapbuf_size64_14_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_15_sram;
wire [0:6] mux_tree_tapbuf_size64_15_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_16_sram;
wire [0:6] mux_tree_tapbuf_size64_16_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_17_sram;
wire [0:6] mux_tree_tapbuf_size64_17_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_18_sram;
wire [0:6] mux_tree_tapbuf_size64_18_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_19_sram;
wire [0:6] mux_tree_tapbuf_size64_19_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_1_sram;
wire [0:6] mux_tree_tapbuf_size64_1_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_20_sram;
wire [0:6] mux_tree_tapbuf_size64_20_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_21_sram;
wire [0:6] mux_tree_tapbuf_size64_21_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_22_sram;
wire [0:6] mux_tree_tapbuf_size64_22_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_23_sram;
wire [0:6] mux_tree_tapbuf_size64_23_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_24_sram;
wire [0:6] mux_tree_tapbuf_size64_24_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_25_sram;
wire [0:6] mux_tree_tapbuf_size64_25_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_26_sram;
wire [0:6] mux_tree_tapbuf_size64_26_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_27_sram;
wire [0:6] mux_tree_tapbuf_size64_27_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_28_sram;
wire [0:6] mux_tree_tapbuf_size64_28_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_29_sram;
wire [0:6] mux_tree_tapbuf_size64_29_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_2_sram;
wire [0:6] mux_tree_tapbuf_size64_2_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_30_sram;
wire [0:6] mux_tree_tapbuf_size64_30_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_31_sram;
wire [0:6] mux_tree_tapbuf_size64_31_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_32_sram;
wire [0:6] mux_tree_tapbuf_size64_32_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_33_sram;
wire [0:6] mux_tree_tapbuf_size64_33_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_34_sram;
wire [0:6] mux_tree_tapbuf_size64_34_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_35_sram;
wire [0:6] mux_tree_tapbuf_size64_35_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_36_sram;
wire [0:6] mux_tree_tapbuf_size64_36_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_37_sram;
wire [0:6] mux_tree_tapbuf_size64_37_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_38_sram;
wire [0:6] mux_tree_tapbuf_size64_38_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_39_sram;
wire [0:6] mux_tree_tapbuf_size64_39_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_3_sram;
wire [0:6] mux_tree_tapbuf_size64_3_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_40_sram;
wire [0:6] mux_tree_tapbuf_size64_40_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_41_sram;
wire [0:6] mux_tree_tapbuf_size64_41_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_42_sram;
wire [0:6] mux_tree_tapbuf_size64_42_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_43_sram;
wire [0:6] mux_tree_tapbuf_size64_43_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_44_sram;
wire [0:6] mux_tree_tapbuf_size64_44_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_45_sram;
wire [0:6] mux_tree_tapbuf_size64_45_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_46_sram;
wire [0:6] mux_tree_tapbuf_size64_46_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_47_sram;
wire [0:6] mux_tree_tapbuf_size64_47_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_48_sram;
wire [0:6] mux_tree_tapbuf_size64_48_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_49_sram;
wire [0:6] mux_tree_tapbuf_size64_49_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_4_sram;
wire [0:6] mux_tree_tapbuf_size64_4_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_50_sram;
wire [0:6] mux_tree_tapbuf_size64_50_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_51_sram;
wire [0:6] mux_tree_tapbuf_size64_51_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_52_sram;
wire [0:6] mux_tree_tapbuf_size64_52_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_53_sram;
wire [0:6] mux_tree_tapbuf_size64_53_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_54_sram;
wire [0:6] mux_tree_tapbuf_size64_54_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_55_sram;
wire [0:6] mux_tree_tapbuf_size64_55_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_56_sram;
wire [0:6] mux_tree_tapbuf_size64_56_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_57_sram;
wire [0:6] mux_tree_tapbuf_size64_57_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_58_sram;
wire [0:6] mux_tree_tapbuf_size64_58_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_59_sram;
wire [0:6] mux_tree_tapbuf_size64_59_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_5_sram;
wire [0:6] mux_tree_tapbuf_size64_5_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_60_sram;
wire [0:6] mux_tree_tapbuf_size64_60_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_61_sram;
wire [0:6] mux_tree_tapbuf_size64_61_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_62_sram;
wire [0:6] mux_tree_tapbuf_size64_62_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_63_sram;
wire [0:6] mux_tree_tapbuf_size64_63_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_64_sram;
wire [0:6] mux_tree_tapbuf_size64_64_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_65_sram;
wire [0:6] mux_tree_tapbuf_size64_65_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_66_sram;
wire [0:6] mux_tree_tapbuf_size64_66_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_67_sram;
wire [0:6] mux_tree_tapbuf_size64_67_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_68_sram;
wire [0:6] mux_tree_tapbuf_size64_68_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_69_sram;
wire [0:6] mux_tree_tapbuf_size64_69_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_6_sram;
wire [0:6] mux_tree_tapbuf_size64_6_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_70_sram;
wire [0:6] mux_tree_tapbuf_size64_70_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_71_sram;
wire [0:6] mux_tree_tapbuf_size64_71_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_72_sram;
wire [0:6] mux_tree_tapbuf_size64_72_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_73_sram;
wire [0:6] mux_tree_tapbuf_size64_73_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_74_sram;
wire [0:6] mux_tree_tapbuf_size64_74_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_75_sram;
wire [0:6] mux_tree_tapbuf_size64_75_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_76_sram;
wire [0:6] mux_tree_tapbuf_size64_76_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_77_sram;
wire [0:6] mux_tree_tapbuf_size64_77_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_78_sram;
wire [0:6] mux_tree_tapbuf_size64_78_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_79_sram;
wire [0:6] mux_tree_tapbuf_size64_79_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_7_sram;
wire [0:6] mux_tree_tapbuf_size64_7_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_80_sram;
wire [0:6] mux_tree_tapbuf_size64_80_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_81_sram;
wire [0:6] mux_tree_tapbuf_size64_81_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_82_sram;
wire [0:6] mux_tree_tapbuf_size64_82_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_83_sram;
wire [0:6] mux_tree_tapbuf_size64_83_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_84_sram;
wire [0:6] mux_tree_tapbuf_size64_84_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_85_sram;
wire [0:6] mux_tree_tapbuf_size64_85_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_86_sram;
wire [0:6] mux_tree_tapbuf_size64_86_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_87_sram;
wire [0:6] mux_tree_tapbuf_size64_87_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_88_sram;
wire [0:6] mux_tree_tapbuf_size64_88_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_89_sram;
wire [0:6] mux_tree_tapbuf_size64_89_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_8_sram;
wire [0:6] mux_tree_tapbuf_size64_8_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_90_sram;
wire [0:6] mux_tree_tapbuf_size64_90_sram_inv;
wire [0:6] mux_tree_tapbuf_size64_9_sram;
wire [0:6] mux_tree_tapbuf_size64_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size64_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size64_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[0] = chany_bottom_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[2];
// ----- Local connection due to Wire 3 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[3];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[4] = chany_bottom_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[6];
// ----- Local connection due to Wire 7 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[7];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[8] = chany_bottom_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[10];
// ----- Local connection due to Wire 11 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[11];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[12] = chany_bottom_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[14];
// ----- Local connection due to Wire 15 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[15];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[16] = chany_bottom_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[18];
// ----- Local connection due to Wire 19 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[19];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[20] = chany_bottom_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[22];
// ----- Local connection due to Wire 23 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[23];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[24] = chany_bottom_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[26];
// ----- Local connection due to Wire 27 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[27];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[28] = chany_bottom_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[30];
// ----- Local connection due to Wire 31 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[31];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[32] = chany_bottom_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[34];
// ----- Local connection due to Wire 35 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[35];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[36] = chany_bottom_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[38];
// ----- Local connection due to Wire 39 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[39];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[40] = chany_bottom_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[42];
// ----- Local connection due to Wire 43 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[43];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[44] = chany_bottom_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[46];
// ----- Local connection due to Wire 47 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[47];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[48] = chany_bottom_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[50];
// ----- Local connection due to Wire 51 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[51];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[52] = chany_bottom_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[54];
// ----- Local connection due to Wire 55 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[55];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[56] = chany_bottom_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[58];
// ----- Local connection due to Wire 59 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[59];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[60] = chany_bottom_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[62];
// ----- Local connection due to Wire 63 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[63];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[64] = chany_bottom_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[66];
// ----- Local connection due to Wire 67 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[67];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[68] = chany_bottom_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[70];
// ----- Local connection due to Wire 71 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[71];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[72] = chany_bottom_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[74];
// ----- Local connection due to Wire 75 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[75];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[76] = chany_bottom_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[78];
// ----- Local connection due to Wire 79 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[79];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[80] = chany_bottom_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[82];
// ----- Local connection due to Wire 83 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[83];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[84] = chany_bottom_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[86];
// ----- Local connection due to Wire 87 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[87];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[88] = chany_bottom_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[90];
// ----- Local connection due to Wire 91 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[91];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[92] = chany_bottom_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[94];
// ----- Local connection due to Wire 95 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[95];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[96] = chany_bottom_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[98];
// ----- Local connection due to Wire 99 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[99];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[100] = chany_bottom_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[102];
// ----- Local connection due to Wire 103 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[103];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[104] = chany_bottom_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[106];
// ----- Local connection due to Wire 107 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[107];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[108] = chany_bottom_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[110];
// ----- Local connection due to Wire 111 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[111];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[112] = chany_bottom_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[114];
// ----- Local connection due to Wire 115 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[115];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[116] = chany_bottom_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[118];
// ----- Local connection due to Wire 119 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[119];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[120] = chany_bottom_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[122];
// ----- Local connection due to Wire 123 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[123];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[124] = chany_bottom_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[126];
// ----- Local connection due to Wire 127 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[127];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[128] = chany_bottom_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[130];
// ----- Local connection due to Wire 131 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[131];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[132] = chany_bottom_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[134];
// ----- Local connection due to Wire 135 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[135];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[136] = chany_bottom_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[138];
// ----- Local connection due to Wire 139 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[139];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[140] = chany_bottom_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[142];
// ----- Local connection due to Wire 143 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[143];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[144] = chany_bottom_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[146];
// ----- Local connection due to Wire 147 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[147];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[148] = chany_bottom_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[150];
// ----- Local connection due to Wire 151 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[151];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[152] = chany_bottom_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[154];
// ----- Local connection due to Wire 155 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[155];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[156] = chany_bottom_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[158];
// ----- Local connection due to Wire 159 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[159];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[160] = chany_bottom_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[162];
// ----- Local connection due to Wire 163 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[163];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[164] = chany_bottom_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[166];
// ----- Local connection due to Wire 167 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[167];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[168] = chany_bottom_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[170];
// ----- Local connection due to Wire 171 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[171];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[172] = chany_bottom_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[174];
// ----- Local connection due to Wire 175 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[175];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[176] = chany_bottom_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[178];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[179];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[180] = chany_bottom_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[182];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[183];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[184] = chany_bottom_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[186];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[187];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[188] = chany_bottom_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[0] = chany_top_in[0];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[1];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[2];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[3];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[4] = chany_top_in[4];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[5];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[6];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[7];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[8] = chany_top_in[8];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[9];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[10];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[11];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[12] = chany_top_in[12];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[13];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[14];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[15];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[16] = chany_top_in[16];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[17];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[18];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[19];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[20] = chany_top_in[20];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[21];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[22];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[23];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[24] = chany_top_in[24];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[25];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[26];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[27];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[28] = chany_top_in[28];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[29];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[30];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[31];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[32] = chany_top_in[32];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[33];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[34];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[35];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[36] = chany_top_in[36];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[37];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[38];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[39];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[40] = chany_top_in[40];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[41];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[42];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[43];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[44] = chany_top_in[44];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[45];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[46];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[47];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[48] = chany_top_in[48];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[49];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[50];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[51];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[52] = chany_top_in[52];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[53];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[54];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[55];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[56] = chany_top_in[56];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[57];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[58];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[59];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[60] = chany_top_in[60];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[61];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[62];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[63];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[64] = chany_top_in[64];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[65];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[66];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[67];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[68] = chany_top_in[68];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[69];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[70];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[71];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[72] = chany_top_in[72];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[73];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[74];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[75];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[76] = chany_top_in[76];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[77];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[78];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[79];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[80] = chany_top_in[80];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[81];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[82];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[83];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[84] = chany_top_in[84];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[85];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[86];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[87];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[88] = chany_top_in[88];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[89];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[90];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[91];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[92] = chany_top_in[92];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[93];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[94];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[95];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[96] = chany_top_in[96];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[97];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[98];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[99];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[100] = chany_top_in[100];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[101];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[102];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[103];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[104] = chany_top_in[104];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[105] = chany_top_in[105];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[106] = chany_top_in[106];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[107] = chany_top_in[107];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[108] = chany_top_in[108];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chany_top_in[109];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[110] = chany_top_in[110];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[111] = chany_top_in[111];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[112] = chany_top_in[112];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[113] = chany_top_in[113];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[114] = chany_top_in[114];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[115] = chany_top_in[115];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[116] = chany_top_in[116];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[117] = chany_top_in[117];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chany_top_in[118];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chany_top_in[119];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[120] = chany_top_in[120];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[121] = chany_top_in[121];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[122] = chany_top_in[122];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[123] = chany_top_in[123];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[124] = chany_top_in[124];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[125] = chany_top_in[125];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[126] = chany_top_in[126];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[127] = chany_top_in[127];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[128] = chany_top_in[128];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chany_top_in[129];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[130] = chany_top_in[130];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[131] = chany_top_in[131];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[132] = chany_top_in[132];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[133] = chany_top_in[133];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[134] = chany_top_in[134];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[135] = chany_top_in[135];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[136] = chany_top_in[136];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[137] = chany_top_in[137];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chany_top_in[138];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chany_top_in[139];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[140] = chany_top_in[140];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[141] = chany_top_in[141];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[142] = chany_top_in[142];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[143] = chany_top_in[143];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[144] = chany_top_in[144];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[145] = chany_top_in[145];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[146] = chany_top_in[146];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[147] = chany_top_in[147];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[148] = chany_top_in[148];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chany_top_in[149];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[150] = chany_top_in[150];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[151] = chany_top_in[151];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[152] = chany_top_in[152];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[153] = chany_top_in[153];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[154] = chany_top_in[154];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[155] = chany_top_in[155];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[156] = chany_top_in[156];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[157] = chany_top_in[157];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[158] = chany_top_in[158];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[159] = chany_top_in[159];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[160] = chany_top_in[160];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[161] = chany_top_in[161];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[162] = chany_top_in[162];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[163] = chany_top_in[163];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[164] = chany_top_in[164];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[165] = chany_top_in[165];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[166] = chany_top_in[166];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[167] = chany_top_in[167];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[168] = chany_top_in[168];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[169] = chany_top_in[169];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[170] = chany_top_in[170];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[171] = chany_top_in[171];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[172] = chany_top_in[172];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[173] = chany_top_in[173];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[174] = chany_top_in[174];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[175] = chany_top_in[175];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[176] = chany_top_in[176];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[177] = chany_top_in[177];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[178] = chany_top_in[178];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[179] = chany_top_in[179];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[180] = chany_top_in[180];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[181] = chany_top_in[181];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[182] = chany_top_in[182];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[183] = chany_top_in[183];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[184] = chany_top_in[184];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[185] = chany_top_in[185];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[186] = chany_top_in[186];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[187] = chany_top_in[187];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[188] = chany_top_in[188];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size64 mux_left_ipin_0 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_0_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_0_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_I_3_));

	mux_tree_tapbuf_size64 mux_left_ipin_1 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_1_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_1_sram_inv[0:6]),
		.out(right_grid_left_width_0_height_0_subtile_0__pin_I_7_));

	mux_tree_tapbuf_size64 mux_right_ipin_0 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_2_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_2_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_));

	mux_tree_tapbuf_size64 mux_right_ipin_1 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_3_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_3_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_));

	mux_tree_tapbuf_size64 mux_right_ipin_2 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_4_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_4_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_));

	mux_tree_tapbuf_size64 mux_right_ipin_3 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_5_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_5_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_));

	mux_tree_tapbuf_size64 mux_right_ipin_4 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_6_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_6_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_));

	mux_tree_tapbuf_size64 mux_right_ipin_5 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_7_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_7_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_));

	mux_tree_tapbuf_size64 mux_right_ipin_6 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_8_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_8_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_));

	mux_tree_tapbuf_size64 mux_right_ipin_7 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_9_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_9_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_));

	mux_tree_tapbuf_size64 mux_right_ipin_8 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_10_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_10_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_));

	mux_tree_tapbuf_size64 mux_right_ipin_9 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_11_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_11_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_));

	mux_tree_tapbuf_size64 mux_right_ipin_10 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_12_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_12_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_));

	mux_tree_tapbuf_size64 mux_right_ipin_11 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_13_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_13_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_));

	mux_tree_tapbuf_size64 mux_right_ipin_12 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_14_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_14_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_));

	mux_tree_tapbuf_size64 mux_right_ipin_13 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_15_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_15_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_));

	mux_tree_tapbuf_size64 mux_right_ipin_14 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_16_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_16_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_));

	mux_tree_tapbuf_size64 mux_right_ipin_15 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_17_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_17_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_));

	mux_tree_tapbuf_size64 mux_right_ipin_16 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_18_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_18_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_));

	mux_tree_tapbuf_size64 mux_right_ipin_17 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_19_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_19_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_));

	mux_tree_tapbuf_size64 mux_right_ipin_18 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_20_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_20_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_));

	mux_tree_tapbuf_size64 mux_right_ipin_19 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_21_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_21_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_));

	mux_tree_tapbuf_size64 mux_right_ipin_20 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_22_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_22_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_));

	mux_tree_tapbuf_size64 mux_right_ipin_21 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_23_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_23_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_));

	mux_tree_tapbuf_size64 mux_right_ipin_22 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_24_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_24_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_));

	mux_tree_tapbuf_size64 mux_right_ipin_23 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_25_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_25_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_));

	mux_tree_tapbuf_size64 mux_right_ipin_24 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_26_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_26_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_));

	mux_tree_tapbuf_size64 mux_right_ipin_25 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_27_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_27_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_));

	mux_tree_tapbuf_size64 mux_right_ipin_26 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_28_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_28_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_));

	mux_tree_tapbuf_size64 mux_right_ipin_27 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_29_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_29_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_));

	mux_tree_tapbuf_size64 mux_right_ipin_28 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_30_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_30_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_));

	mux_tree_tapbuf_size64 mux_right_ipin_29 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_31_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_31_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_));

	mux_tree_tapbuf_size64 mux_right_ipin_30 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_32_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_32_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_));

	mux_tree_tapbuf_size64 mux_right_ipin_31 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_33_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_33_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_));

	mux_tree_tapbuf_size64 mux_right_ipin_32 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_34_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_34_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_));

	mux_tree_tapbuf_size64 mux_right_ipin_33 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_35_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_35_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_));

	mux_tree_tapbuf_size64 mux_right_ipin_34 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_36_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_36_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_));

	mux_tree_tapbuf_size64 mux_right_ipin_35 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_37_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_37_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_));

	mux_tree_tapbuf_size64 mux_right_ipin_36 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_38_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_38_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_));

	mux_tree_tapbuf_size64 mux_right_ipin_37 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_39_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_39_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_));

	mux_tree_tapbuf_size64 mux_right_ipin_38 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_40_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_40_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_));

	mux_tree_tapbuf_size64 mux_right_ipin_39 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_41_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_41_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_));

	mux_tree_tapbuf_size64 mux_right_ipin_40 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_42_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_42_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_));

	mux_tree_tapbuf_size64 mux_right_ipin_41 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_43_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_43_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_));

	mux_tree_tapbuf_size64 mux_right_ipin_42 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_44_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_44_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_));

	mux_tree_tapbuf_size64 mux_right_ipin_43 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_45_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_45_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_));

	mux_tree_tapbuf_size64 mux_right_ipin_44 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_46_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_46_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_));

	mux_tree_tapbuf_size64 mux_right_ipin_45 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_47_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_47_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_));

	mux_tree_tapbuf_size64 mux_right_ipin_46 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_48_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_48_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_));

	mux_tree_tapbuf_size64 mux_right_ipin_47 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_49_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_49_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_));

	mux_tree_tapbuf_size64 mux_right_ipin_48 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_50_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_50_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_));

	mux_tree_tapbuf_size64 mux_right_ipin_49 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_51_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_51_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_));

	mux_tree_tapbuf_size64 mux_right_ipin_50 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_52_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_52_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_));

	mux_tree_tapbuf_size64 mux_right_ipin_51 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_53_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_53_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_));

	mux_tree_tapbuf_size64 mux_right_ipin_52 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_54_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_54_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_));

	mux_tree_tapbuf_size64 mux_right_ipin_53 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_55_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_55_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_));

	mux_tree_tapbuf_size64 mux_right_ipin_54 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_56_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_56_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_));

	mux_tree_tapbuf_size64 mux_right_ipin_55 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_57_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_57_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_));

	mux_tree_tapbuf_size64 mux_right_ipin_56 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_58_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_58_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_));

	mux_tree_tapbuf_size64 mux_right_ipin_57 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_59_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_59_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_));

	mux_tree_tapbuf_size64 mux_right_ipin_58 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_60_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_60_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_));

	mux_tree_tapbuf_size64 mux_right_ipin_59 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_61_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_61_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_));

	mux_tree_tapbuf_size64 mux_right_ipin_60 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_62_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_62_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_));

	mux_tree_tapbuf_size64 mux_right_ipin_61 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_63_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_63_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_));

	mux_tree_tapbuf_size64 mux_right_ipin_62 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_64_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_64_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_));

	mux_tree_tapbuf_size64 mux_right_ipin_63 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_65_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_65_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_));

	mux_tree_tapbuf_size64 mux_right_ipin_64 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_66_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_66_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_));

	mux_tree_tapbuf_size64 mux_right_ipin_65 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_67_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_67_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_));

	mux_tree_tapbuf_size64 mux_right_ipin_66 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_68_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_68_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_));

	mux_tree_tapbuf_size64 mux_right_ipin_67 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_69_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_69_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_));

	mux_tree_tapbuf_size64 mux_right_ipin_68 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_70_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_70_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_));

	mux_tree_tapbuf_size64 mux_right_ipin_69 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_71_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_71_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_));

	mux_tree_tapbuf_size64 mux_right_ipin_70 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_72_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_72_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_));

	mux_tree_tapbuf_size64 mux_right_ipin_71 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_73_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_73_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_));

	mux_tree_tapbuf_size64 mux_right_ipin_72 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_74_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_74_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_));

	mux_tree_tapbuf_size64 mux_right_ipin_73 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_75_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_75_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_));

	mux_tree_tapbuf_size64 mux_right_ipin_74 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_76_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_76_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_));

	mux_tree_tapbuf_size64 mux_right_ipin_75 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_77_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_77_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_));

	mux_tree_tapbuf_size64 mux_right_ipin_76 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_78_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_78_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_));

	mux_tree_tapbuf_size64 mux_right_ipin_77 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_79_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_79_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_));

	mux_tree_tapbuf_size64 mux_right_ipin_78 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_80_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_80_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_));

	mux_tree_tapbuf_size64 mux_right_ipin_79 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_81_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_81_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_));

	mux_tree_tapbuf_size64 mux_right_ipin_80 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_82_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_82_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_));

	mux_tree_tapbuf_size64 mux_right_ipin_81 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_83_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_83_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_));

	mux_tree_tapbuf_size64 mux_right_ipin_82 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_84_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_84_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_));

	mux_tree_tapbuf_size64 mux_right_ipin_83 (
		.in({chany_bottom_in[4], chany_top_in[4], chany_bottom_in[10], chany_top_in[10], chany_bottom_in[16], chany_top_in[16], chany_bottom_in[22], chany_top_in[22], chany_bottom_in[28], chany_top_in[28], chany_bottom_in[34], chany_top_in[34], chany_bottom_in[40], chany_top_in[40], chany_bottom_in[46], chany_top_in[46], chany_bottom_in[52], chany_top_in[52], chany_bottom_in[58], chany_top_in[58], chany_bottom_in[64], chany_top_in[64], chany_bottom_in[70], chany_top_in[70], chany_bottom_in[76], chany_top_in[76], chany_bottom_in[82], chany_top_in[82], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[91], chany_top_in[91], chany_bottom_in[97], chany_top_in[97], chany_bottom_in[103], chany_top_in[103], chany_bottom_in[109], chany_top_in[109], chany_bottom_in[115], chany_top_in[115], chany_bottom_in[121], chany_top_in[121], chany_bottom_in[127], chany_top_in[127], chany_bottom_in[133], chany_top_in[133], chany_bottom_in[139], chany_top_in[139], chany_bottom_in[145], chany_top_in[145], chany_bottom_in[151], chany_top_in[151], chany_bottom_in[157], chany_top_in[157], chany_bottom_in[163], chany_top_in[163], chany_bottom_in[169], chany_top_in[169], chany_bottom_in[175], chany_top_in[175], chany_bottom_in[181], chany_top_in[181], chany_bottom_in[187], chany_top_in[187]}),
		.sram(mux_tree_tapbuf_size64_85_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_85_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_));

	mux_tree_tapbuf_size64 mux_right_ipin_84 (
		.in({chany_bottom_in[5], chany_top_in[5], chany_bottom_in[11], chany_top_in[11], chany_bottom_in[17], chany_top_in[17], chany_bottom_in[23], chany_top_in[23], chany_bottom_in[29], chany_top_in[29], chany_bottom_in[35], chany_top_in[35], chany_bottom_in[41], chany_top_in[41], chany_bottom_in[47], chany_top_in[47], chany_bottom_in[53], chany_top_in[53], chany_bottom_in[59], chany_top_in[59], chany_bottom_in[65], chany_top_in[65], chany_bottom_in[71], chany_top_in[71], chany_bottom_in[77], chany_top_in[77], chany_bottom_in[83], chany_top_in[83], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[92], chany_top_in[92], chany_bottom_in[98], chany_top_in[98], chany_bottom_in[104], chany_top_in[104], chany_bottom_in[110], chany_top_in[110], chany_bottom_in[116], chany_top_in[116], chany_bottom_in[122], chany_top_in[122], chany_bottom_in[128], chany_top_in[128], chany_bottom_in[134], chany_top_in[134], chany_bottom_in[140], chany_top_in[140], chany_bottom_in[146], chany_top_in[146], chany_bottom_in[152], chany_top_in[152], chany_bottom_in[158], chany_top_in[158], chany_bottom_in[164], chany_top_in[164], chany_bottom_in[170], chany_top_in[170], chany_bottom_in[176], chany_top_in[176], chany_bottom_in[182], chany_top_in[182], chany_bottom_in[188], chany_top_in[188]}),
		.sram(mux_tree_tapbuf_size64_86_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_86_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_));

	mux_tree_tapbuf_size64 mux_right_ipin_85 (
		.in({chany_bottom_in[0], chany_top_in[0], chany_bottom_in[6], chany_top_in[6], chany_bottom_in[12], chany_top_in[12], chany_bottom_in[18], chany_top_in[18], chany_bottom_in[24], chany_top_in[24], chany_bottom_in[30], chany_top_in[30], chany_bottom_in[36], chany_top_in[36], chany_bottom_in[42], chany_top_in[42], chany_bottom_in[48], chany_top_in[48], chany_bottom_in[54], chany_top_in[54], chany_bottom_in[60], chany_top_in[60], chany_bottom_in[66], chany_top_in[66], chany_bottom_in[72], chany_top_in[72], chany_bottom_in[78], chany_top_in[78], chany_bottom_in[84], chany_top_in[84], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[93], chany_top_in[93], chany_bottom_in[99], chany_top_in[99], chany_bottom_in[105], chany_top_in[105], chany_bottom_in[111], chany_top_in[111], chany_bottom_in[117], chany_top_in[117], chany_bottom_in[123], chany_top_in[123], chany_bottom_in[129], chany_top_in[129], chany_bottom_in[135], chany_top_in[135], chany_bottom_in[141], chany_top_in[141], chany_bottom_in[147], chany_top_in[147], chany_bottom_in[153], chany_top_in[153], chany_bottom_in[159], chany_top_in[159], chany_bottom_in[165], chany_top_in[165], chany_bottom_in[171], chany_top_in[171], chany_bottom_in[177], chany_top_in[177], chany_bottom_in[183], chany_top_in[183]}),
		.sram(mux_tree_tapbuf_size64_87_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_87_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_));

	mux_tree_tapbuf_size64 mux_right_ipin_86 (
		.in({chany_bottom_in[1], chany_top_in[1], chany_bottom_in[7], chany_top_in[7], chany_bottom_in[13], chany_top_in[13], chany_bottom_in[19], chany_top_in[19], chany_bottom_in[25], chany_top_in[25], chany_bottom_in[31], chany_top_in[31], chany_bottom_in[37], chany_top_in[37], chany_bottom_in[43], chany_top_in[43], chany_bottom_in[49], chany_top_in[49], chany_bottom_in[55], chany_top_in[55], chany_bottom_in[61], chany_top_in[61], chany_bottom_in[67], chany_top_in[67], chany_bottom_in[73], chany_top_in[73], chany_bottom_in[79], chany_top_in[79], chany_bottom_in[85], chany_top_in[85], chany_bottom_in[88], chany_top_in[88], chany_bottom_in[94], chany_top_in[94], chany_bottom_in[100], chany_top_in[100], chany_bottom_in[106], chany_top_in[106], chany_bottom_in[112], chany_top_in[112], chany_bottom_in[118], chany_top_in[118], chany_bottom_in[124], chany_top_in[124], chany_bottom_in[130], chany_top_in[130], chany_bottom_in[136], chany_top_in[136], chany_bottom_in[142], chany_top_in[142], chany_bottom_in[148], chany_top_in[148], chany_bottom_in[154], chany_top_in[154], chany_bottom_in[160], chany_top_in[160], chany_bottom_in[166], chany_top_in[166], chany_bottom_in[172], chany_top_in[172], chany_bottom_in[178], chany_top_in[178], chany_bottom_in[184], chany_top_in[184]}),
		.sram(mux_tree_tapbuf_size64_88_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_88_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_));

	mux_tree_tapbuf_size64 mux_right_ipin_87 (
		.in({chany_bottom_in[2], chany_top_in[2], chany_bottom_in[8], chany_top_in[8], chany_bottom_in[14], chany_top_in[14], chany_bottom_in[20], chany_top_in[20], chany_bottom_in[26], chany_top_in[26], chany_bottom_in[32], chany_top_in[32], chany_bottom_in[38], chany_top_in[38], chany_bottom_in[44], chany_top_in[44], chany_bottom_in[50], chany_top_in[50], chany_bottom_in[56], chany_top_in[56], chany_bottom_in[62], chany_top_in[62], chany_bottom_in[68], chany_top_in[68], chany_bottom_in[74], chany_top_in[74], chany_bottom_in[80], chany_top_in[80], chany_bottom_in[86], chany_top_in[86], chany_bottom_in[89], chany_top_in[89], chany_bottom_in[95], chany_top_in[95], chany_bottom_in[101], chany_top_in[101], chany_bottom_in[107], chany_top_in[107], chany_bottom_in[113], chany_top_in[113], chany_bottom_in[119], chany_top_in[119], chany_bottom_in[125], chany_top_in[125], chany_bottom_in[131], chany_top_in[131], chany_bottom_in[137], chany_top_in[137], chany_bottom_in[143], chany_top_in[143], chany_bottom_in[149], chany_top_in[149], chany_bottom_in[155], chany_top_in[155], chany_bottom_in[161], chany_top_in[161], chany_bottom_in[167], chany_top_in[167], chany_bottom_in[173], chany_top_in[173], chany_bottom_in[179], chany_top_in[179], chany_bottom_in[185], chany_top_in[185]}),
		.sram(mux_tree_tapbuf_size64_89_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_89_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_));

	mux_tree_tapbuf_size64 mux_right_ipin_88 (
		.in({chany_bottom_in[3], chany_top_in[3], chany_bottom_in[9], chany_top_in[9], chany_bottom_in[15], chany_top_in[15], chany_bottom_in[21], chany_top_in[21], chany_bottom_in[27], chany_top_in[27], chany_bottom_in[33], chany_top_in[33], chany_bottom_in[39], chany_top_in[39], chany_bottom_in[45], chany_top_in[45], chany_bottom_in[51], chany_top_in[51], chany_bottom_in[57], chany_top_in[57], chany_bottom_in[63], chany_top_in[63], chany_bottom_in[69], chany_top_in[69], chany_bottom_in[75], chany_top_in[75], chany_bottom_in[81], chany_top_in[81], chany_bottom_in[87], chany_top_in[87], chany_bottom_in[90], chany_top_in[90], chany_bottom_in[96], chany_top_in[96], chany_bottom_in[102], chany_top_in[102], chany_bottom_in[108], chany_top_in[108], chany_bottom_in[114], chany_top_in[114], chany_bottom_in[120], chany_top_in[120], chany_bottom_in[126], chany_top_in[126], chany_bottom_in[132], chany_top_in[132], chany_bottom_in[138], chany_top_in[138], chany_bottom_in[144], chany_top_in[144], chany_bottom_in[150], chany_top_in[150], chany_bottom_in[156], chany_top_in[156], chany_bottom_in[162], chany_top_in[162], chany_bottom_in[168], chany_top_in[168], chany_bottom_in[174], chany_top_in[174], chany_bottom_in[180], chany_top_in[180], chany_bottom_in[186], chany_top_in[186]}),
		.sram(mux_tree_tapbuf_size64_90_sram[0:6]),
		.sram_inv(mux_tree_tapbuf_size64_90_sram_inv[0:6]),
		.out(left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_));

	mux_tree_tapbuf_size64_mem mem_left_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size64_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_0_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_0_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_left_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_1_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_1_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_2_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_2_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_3_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_3_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_4_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_4_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_5_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_5_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_6_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_6_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_7_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_7_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_8_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_8_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_9_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_9_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_10_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_10_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_11_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_11_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_12_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_12_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_13_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_13_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_14_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_14_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_15_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_15_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_16_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_16_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_17_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_17_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_18_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_18_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_19_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_19_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_20_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_20_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_21_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_21_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_22_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_22_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_23_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_23_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_24_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_24_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_25_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_25_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_26_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_26_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_27_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_27_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_28_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_28_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_29_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_29_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_30_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_30_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_31_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_31_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_32_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_32_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_33_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_33_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_34_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_34_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_35_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_35_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_36_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_36_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_37_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_37_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_38_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_38_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_39_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_39_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_40_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_40_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_41_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_41_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_42_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_42_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_43_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_43_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_44_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_44_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_45_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_45_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_46_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_46_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_47_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_47_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_48_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_48_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_49_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_49_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_50_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_50_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_51_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_51_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_52_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_52_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_53_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_53_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_54_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_54_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_55_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_55_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_56_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_56_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_57_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_57_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_58_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_58_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_59_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_59_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_60_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_60_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_61_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_61_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_62_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_62_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_63_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_63_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_64_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_64_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_65_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_65_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_66_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_66_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_67_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_67_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_68_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_68_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_69_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_69_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_70_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_70_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_71_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_71_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_72_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_72_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_73_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_73_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_74_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_74_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_75_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_75_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_76_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_76_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_77_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_77_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_78_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_78_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_79_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_79_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_80_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_80_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_81_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_81_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_82_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_82_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_83_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_83_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_84_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_84_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_85_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_85_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_86_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_86_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_87_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_87_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_88_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_88_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size64_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_89_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_89_sram_inv[0:6]));

	mux_tree_tapbuf_size64_mem mem_right_ipin_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size64_mem_89_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size64_90_sram[0:6]),
		.mem_outb(mux_tree_tapbuf_size64_90_sram_inv[0:6]));

endmodule
// ----- END Verilog module for cby_1__2_ -----

//----- Default net type -----
`default_nettype wire




