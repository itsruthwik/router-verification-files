//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][4]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul  7 20:54:34 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__4_ -----
module sb_0__4_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:295] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:295] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:295] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:295] chany_top_out;
//----- OUTPUT PORTS -----
output [0:295] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:295] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_100_sram;
wire [0:1] mux_tree_tapbuf_size3_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_101_sram;
wire [0:1] mux_tree_tapbuf_size3_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_102_sram;
wire [0:1] mux_tree_tapbuf_size3_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_103_sram;
wire [0:1] mux_tree_tapbuf_size3_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_104_sram;
wire [0:1] mux_tree_tapbuf_size3_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_105_sram;
wire [0:1] mux_tree_tapbuf_size3_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_106_sram;
wire [0:1] mux_tree_tapbuf_size3_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_107_sram;
wire [0:1] mux_tree_tapbuf_size3_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_108_sram;
wire [0:1] mux_tree_tapbuf_size3_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_109_sram;
wire [0:1] mux_tree_tapbuf_size3_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_110_sram;
wire [0:1] mux_tree_tapbuf_size3_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_111_sram;
wire [0:1] mux_tree_tapbuf_size3_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_112_sram;
wire [0:1] mux_tree_tapbuf_size3_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_113_sram;
wire [0:1] mux_tree_tapbuf_size3_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_114_sram;
wire [0:1] mux_tree_tapbuf_size3_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_115_sram;
wire [0:1] mux_tree_tapbuf_size3_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_116_sram;
wire [0:1] mux_tree_tapbuf_size3_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_117_sram;
wire [0:1] mux_tree_tapbuf_size3_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_118_sram;
wire [0:1] mux_tree_tapbuf_size3_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_119_sram;
wire [0:1] mux_tree_tapbuf_size3_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_120_sram;
wire [0:1] mux_tree_tapbuf_size3_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_121_sram;
wire [0:1] mux_tree_tapbuf_size3_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_122_sram;
wire [0:1] mux_tree_tapbuf_size3_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_123_sram;
wire [0:1] mux_tree_tapbuf_size3_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_124_sram;
wire [0:1] mux_tree_tapbuf_size3_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_125_sram;
wire [0:1] mux_tree_tapbuf_size3_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_126_sram;
wire [0:1] mux_tree_tapbuf_size3_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_127_sram;
wire [0:1] mux_tree_tapbuf_size3_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_128_sram;
wire [0:1] mux_tree_tapbuf_size3_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_129_sram;
wire [0:1] mux_tree_tapbuf_size3_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_130_sram;
wire [0:1] mux_tree_tapbuf_size3_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_131_sram;
wire [0:1] mux_tree_tapbuf_size3_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_132_sram;
wire [0:1] mux_tree_tapbuf_size3_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_133_sram;
wire [0:1] mux_tree_tapbuf_size3_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_134_sram;
wire [0:1] mux_tree_tapbuf_size3_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_135_sram;
wire [0:1] mux_tree_tapbuf_size3_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_136_sram;
wire [0:1] mux_tree_tapbuf_size3_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_137_sram;
wire [0:1] mux_tree_tapbuf_size3_137_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_138_sram;
wire [0:1] mux_tree_tapbuf_size3_138_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_139_sram;
wire [0:1] mux_tree_tapbuf_size3_139_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_140_sram;
wire [0:1] mux_tree_tapbuf_size3_140_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_141_sram;
wire [0:1] mux_tree_tapbuf_size3_141_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_142_sram;
wire [0:1] mux_tree_tapbuf_size3_142_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_143_sram;
wire [0:1] mux_tree_tapbuf_size3_143_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_144_sram;
wire [0:1] mux_tree_tapbuf_size3_144_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_145_sram;
wire [0:1] mux_tree_tapbuf_size3_145_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_146_sram;
wire [0:1] mux_tree_tapbuf_size3_146_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_147_sram;
wire [0:1] mux_tree_tapbuf_size3_147_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_148_sram;
wire [0:1] mux_tree_tapbuf_size3_148_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_149_sram;
wire [0:1] mux_tree_tapbuf_size3_149_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_150_sram;
wire [0:1] mux_tree_tapbuf_size3_150_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_151_sram;
wire [0:1] mux_tree_tapbuf_size3_151_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_152_sram;
wire [0:1] mux_tree_tapbuf_size3_152_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_153_sram;
wire [0:1] mux_tree_tapbuf_size3_153_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_154_sram;
wire [0:1] mux_tree_tapbuf_size3_154_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_155_sram;
wire [0:1] mux_tree_tapbuf_size3_155_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_156_sram;
wire [0:1] mux_tree_tapbuf_size3_156_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_157_sram;
wire [0:1] mux_tree_tapbuf_size3_157_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_158_sram;
wire [0:1] mux_tree_tapbuf_size3_158_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_159_sram;
wire [0:1] mux_tree_tapbuf_size3_159_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_160_sram;
wire [0:1] mux_tree_tapbuf_size3_160_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_161_sram;
wire [0:1] mux_tree_tapbuf_size3_161_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_162_sram;
wire [0:1] mux_tree_tapbuf_size3_162_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_163_sram;
wire [0:1] mux_tree_tapbuf_size3_163_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_164_sram;
wire [0:1] mux_tree_tapbuf_size3_164_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_165_sram;
wire [0:1] mux_tree_tapbuf_size3_165_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_166_sram;
wire [0:1] mux_tree_tapbuf_size3_166_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_167_sram;
wire [0:1] mux_tree_tapbuf_size3_167_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_168_sram;
wire [0:1] mux_tree_tapbuf_size3_168_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_169_sram;
wire [0:1] mux_tree_tapbuf_size3_169_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_170_sram;
wire [0:1] mux_tree_tapbuf_size3_170_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_171_sram;
wire [0:1] mux_tree_tapbuf_size3_171_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_172_sram;
wire [0:1] mux_tree_tapbuf_size3_172_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_173_sram;
wire [0:1] mux_tree_tapbuf_size3_173_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_174_sram;
wire [0:1] mux_tree_tapbuf_size3_174_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_175_sram;
wire [0:1] mux_tree_tapbuf_size3_175_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_176_sram;
wire [0:1] mux_tree_tapbuf_size3_176_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_177_sram;
wire [0:1] mux_tree_tapbuf_size3_177_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_178_sram;
wire [0:1] mux_tree_tapbuf_size3_178_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_179_sram;
wire [0:1] mux_tree_tapbuf_size3_179_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_180_sram;
wire [0:1] mux_tree_tapbuf_size3_180_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_181_sram;
wire [0:1] mux_tree_tapbuf_size3_181_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_182_sram;
wire [0:1] mux_tree_tapbuf_size3_182_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_183_sram;
wire [0:1] mux_tree_tapbuf_size3_183_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_184_sram;
wire [0:1] mux_tree_tapbuf_size3_184_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_185_sram;
wire [0:1] mux_tree_tapbuf_size3_185_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_186_sram;
wire [0:1] mux_tree_tapbuf_size3_186_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_187_sram;
wire [0:1] mux_tree_tapbuf_size3_187_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_188_sram;
wire [0:1] mux_tree_tapbuf_size3_188_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_189_sram;
wire [0:1] mux_tree_tapbuf_size3_189_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_190_sram;
wire [0:1] mux_tree_tapbuf_size3_190_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_191_sram;
wire [0:1] mux_tree_tapbuf_size3_191_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_192_sram;
wire [0:1] mux_tree_tapbuf_size3_192_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_193_sram;
wire [0:1] mux_tree_tapbuf_size3_193_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_194_sram;
wire [0:1] mux_tree_tapbuf_size3_194_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_195_sram;
wire [0:1] mux_tree_tapbuf_size3_195_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_196_sram;
wire [0:1] mux_tree_tapbuf_size3_196_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_197_sram;
wire [0:1] mux_tree_tapbuf_size3_197_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_198_sram;
wire [0:1] mux_tree_tapbuf_size3_198_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_199_sram;
wire [0:1] mux_tree_tapbuf_size3_199_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_200_sram;
wire [0:1] mux_tree_tapbuf_size3_200_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_201_sram;
wire [0:1] mux_tree_tapbuf_size3_201_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_202_sram;
wire [0:1] mux_tree_tapbuf_size3_202_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_203_sram;
wire [0:1] mux_tree_tapbuf_size3_203_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_204_sram;
wire [0:1] mux_tree_tapbuf_size3_204_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_205_sram;
wire [0:1] mux_tree_tapbuf_size3_205_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_206_sram;
wire [0:1] mux_tree_tapbuf_size3_206_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_207_sram;
wire [0:1] mux_tree_tapbuf_size3_207_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_208_sram;
wire [0:1] mux_tree_tapbuf_size3_208_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_209_sram;
wire [0:1] mux_tree_tapbuf_size3_209_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_210_sram;
wire [0:1] mux_tree_tapbuf_size3_210_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_211_sram;
wire [0:1] mux_tree_tapbuf_size3_211_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_212_sram;
wire [0:1] mux_tree_tapbuf_size3_212_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_213_sram;
wire [0:1] mux_tree_tapbuf_size3_213_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_214_sram;
wire [0:1] mux_tree_tapbuf_size3_214_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_215_sram;
wire [0:1] mux_tree_tapbuf_size3_215_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_216_sram;
wire [0:1] mux_tree_tapbuf_size3_216_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_217_sram;
wire [0:1] mux_tree_tapbuf_size3_217_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_218_sram;
wire [0:1] mux_tree_tapbuf_size3_218_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_219_sram;
wire [0:1] mux_tree_tapbuf_size3_219_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_220_sram;
wire [0:1] mux_tree_tapbuf_size3_220_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_221_sram;
wire [0:1] mux_tree_tapbuf_size3_221_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_222_sram;
wire [0:1] mux_tree_tapbuf_size3_222_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_223_sram;
wire [0:1] mux_tree_tapbuf_size3_223_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_224_sram;
wire [0:1] mux_tree_tapbuf_size3_224_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_225_sram;
wire [0:1] mux_tree_tapbuf_size3_225_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_226_sram;
wire [0:1] mux_tree_tapbuf_size3_226_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_227_sram;
wire [0:1] mux_tree_tapbuf_size3_227_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_228_sram;
wire [0:1] mux_tree_tapbuf_size3_228_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_229_sram;
wire [0:1] mux_tree_tapbuf_size3_229_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_230_sram;
wire [0:1] mux_tree_tapbuf_size3_230_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_231_sram;
wire [0:1] mux_tree_tapbuf_size3_231_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_232_sram;
wire [0:1] mux_tree_tapbuf_size3_232_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_233_sram;
wire [0:1] mux_tree_tapbuf_size3_233_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_234_sram;
wire [0:1] mux_tree_tapbuf_size3_234_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_235_sram;
wire [0:1] mux_tree_tapbuf_size3_235_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_236_sram;
wire [0:1] mux_tree_tapbuf_size3_236_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_237_sram;
wire [0:1] mux_tree_tapbuf_size3_237_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_238_sram;
wire [0:1] mux_tree_tapbuf_size3_238_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_239_sram;
wire [0:1] mux_tree_tapbuf_size3_239_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_240_sram;
wire [0:1] mux_tree_tapbuf_size3_240_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_241_sram;
wire [0:1] mux_tree_tapbuf_size3_241_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_242_sram;
wire [0:1] mux_tree_tapbuf_size3_242_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_243_sram;
wire [0:1] mux_tree_tapbuf_size3_243_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_244_sram;
wire [0:1] mux_tree_tapbuf_size3_244_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_245_sram;
wire [0:1] mux_tree_tapbuf_size3_245_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_246_sram;
wire [0:1] mux_tree_tapbuf_size3_246_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_247_sram;
wire [0:1] mux_tree_tapbuf_size3_247_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_248_sram;
wire [0:1] mux_tree_tapbuf_size3_248_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_249_sram;
wire [0:1] mux_tree_tapbuf_size3_249_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_250_sram;
wire [0:1] mux_tree_tapbuf_size3_250_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_251_sram;
wire [0:1] mux_tree_tapbuf_size3_251_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_252_sram;
wire [0:1] mux_tree_tapbuf_size3_252_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_253_sram;
wire [0:1] mux_tree_tapbuf_size3_253_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_254_sram;
wire [0:1] mux_tree_tapbuf_size3_254_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_255_sram;
wire [0:1] mux_tree_tapbuf_size3_255_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_256_sram;
wire [0:1] mux_tree_tapbuf_size3_256_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_257_sram;
wire [0:1] mux_tree_tapbuf_size3_257_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_258_sram;
wire [0:1] mux_tree_tapbuf_size3_258_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_259_sram;
wire [0:1] mux_tree_tapbuf_size3_259_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_260_sram;
wire [0:1] mux_tree_tapbuf_size3_260_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_261_sram;
wire [0:1] mux_tree_tapbuf_size3_261_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_262_sram;
wire [0:1] mux_tree_tapbuf_size3_262_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_263_sram;
wire [0:1] mux_tree_tapbuf_size3_263_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_264_sram;
wire [0:1] mux_tree_tapbuf_size3_264_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_265_sram;
wire [0:1] mux_tree_tapbuf_size3_265_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_266_sram;
wire [0:1] mux_tree_tapbuf_size3_266_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_267_sram;
wire [0:1] mux_tree_tapbuf_size3_267_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_268_sram;
wire [0:1] mux_tree_tapbuf_size3_268_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_269_sram;
wire [0:1] mux_tree_tapbuf_size3_269_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_270_sram;
wire [0:1] mux_tree_tapbuf_size3_270_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_271_sram;
wire [0:1] mux_tree_tapbuf_size3_271_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_272_sram;
wire [0:1] mux_tree_tapbuf_size3_272_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_273_sram;
wire [0:1] mux_tree_tapbuf_size3_273_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_274_sram;
wire [0:1] mux_tree_tapbuf_size3_274_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_275_sram;
wire [0:1] mux_tree_tapbuf_size3_275_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_276_sram;
wire [0:1] mux_tree_tapbuf_size3_276_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_277_sram;
wire [0:1] mux_tree_tapbuf_size3_277_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_278_sram;
wire [0:1] mux_tree_tapbuf_size3_278_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_279_sram;
wire [0:1] mux_tree_tapbuf_size3_279_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_280_sram;
wire [0:1] mux_tree_tapbuf_size3_280_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_281_sram;
wire [0:1] mux_tree_tapbuf_size3_281_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_282_sram;
wire [0:1] mux_tree_tapbuf_size3_282_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_283_sram;
wire [0:1] mux_tree_tapbuf_size3_283_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_284_sram;
wire [0:1] mux_tree_tapbuf_size3_284_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_285_sram;
wire [0:1] mux_tree_tapbuf_size3_285_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_286_sram;
wire [0:1] mux_tree_tapbuf_size3_286_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_287_sram;
wire [0:1] mux_tree_tapbuf_size3_287_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_288_sram;
wire [0:1] mux_tree_tapbuf_size3_288_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_289_sram;
wire [0:1] mux_tree_tapbuf_size3_289_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_60_sram;
wire [0:1] mux_tree_tapbuf_size3_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_61_sram;
wire [0:1] mux_tree_tapbuf_size3_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_62_sram;
wire [0:1] mux_tree_tapbuf_size3_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_63_sram;
wire [0:1] mux_tree_tapbuf_size3_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_64_sram;
wire [0:1] mux_tree_tapbuf_size3_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_65_sram;
wire [0:1] mux_tree_tapbuf_size3_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_66_sram;
wire [0:1] mux_tree_tapbuf_size3_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_67_sram;
wire [0:1] mux_tree_tapbuf_size3_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_68_sram;
wire [0:1] mux_tree_tapbuf_size3_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_69_sram;
wire [0:1] mux_tree_tapbuf_size3_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_70_sram;
wire [0:1] mux_tree_tapbuf_size3_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_71_sram;
wire [0:1] mux_tree_tapbuf_size3_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_72_sram;
wire [0:1] mux_tree_tapbuf_size3_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_73_sram;
wire [0:1] mux_tree_tapbuf_size3_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_74_sram;
wire [0:1] mux_tree_tapbuf_size3_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_75_sram;
wire [0:1] mux_tree_tapbuf_size3_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_76_sram;
wire [0:1] mux_tree_tapbuf_size3_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_77_sram;
wire [0:1] mux_tree_tapbuf_size3_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_78_sram;
wire [0:1] mux_tree_tapbuf_size3_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_79_sram;
wire [0:1] mux_tree_tapbuf_size3_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_80_sram;
wire [0:1] mux_tree_tapbuf_size3_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_81_sram;
wire [0:1] mux_tree_tapbuf_size3_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_82_sram;
wire [0:1] mux_tree_tapbuf_size3_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_83_sram;
wire [0:1] mux_tree_tapbuf_size3_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_84_sram;
wire [0:1] mux_tree_tapbuf_size3_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_85_sram;
wire [0:1] mux_tree_tapbuf_size3_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_86_sram;
wire [0:1] mux_tree_tapbuf_size3_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_87_sram;
wire [0:1] mux_tree_tapbuf_size3_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_88_sram;
wire [0:1] mux_tree_tapbuf_size3_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_89_sram;
wire [0:1] mux_tree_tapbuf_size3_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_90_sram;
wire [0:1] mux_tree_tapbuf_size3_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_91_sram;
wire [0:1] mux_tree_tapbuf_size3_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_92_sram;
wire [0:1] mux_tree_tapbuf_size3_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_93_sram;
wire [0:1] mux_tree_tapbuf_size3_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_94_sram;
wire [0:1] mux_tree_tapbuf_size3_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_95_sram;
wire [0:1] mux_tree_tapbuf_size3_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_96_sram;
wire [0:1] mux_tree_tapbuf_size3_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_97_sram;
wire [0:1] mux_tree_tapbuf_size3_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_98_sram;
wire [0:1] mux_tree_tapbuf_size3_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_99_sram;
wire [0:1] mux_tree_tapbuf_size3_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_225_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_226_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_227_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_228_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_229_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_230_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_231_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_232_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_233_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_234_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_235_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_236_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_237_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_238_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_239_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_240_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_241_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_242_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_243_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_244_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_245_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_246_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_247_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_248_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_249_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_250_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_251_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_252_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_253_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_254_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_255_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_256_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_257_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_258_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_259_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_260_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_261_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_262_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_263_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_264_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_265_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_266_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_267_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_268_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_269_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_270_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_271_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_272_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_273_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_274_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_275_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_276_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_277_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_278_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_279_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_280_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_281_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_282_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_283_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_284_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_285_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_286_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_287_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_288_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_289_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_34_sram;
wire [0:2] mux_tree_tapbuf_size5_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_35_sram;
wire [0:2] mux_tree_tapbuf_size5_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_36_sram;
wire [0:2] mux_tree_tapbuf_size5_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_37_sram;
wire [0:2] mux_tree_tapbuf_size5_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_38_sram;
wire [0:2] mux_tree_tapbuf_size5_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_39_sram;
wire [0:2] mux_tree_tapbuf_size5_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_40_sram;
wire [0:2] mux_tree_tapbuf_size5_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_41_sram;
wire [0:2] mux_tree_tapbuf_size5_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_42_sram;
wire [0:2] mux_tree_tapbuf_size5_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_43_sram;
wire [0:2] mux_tree_tapbuf_size5_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_44_sram;
wire [0:2] mux_tree_tapbuf_size5_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_45_sram;
wire [0:2] mux_tree_tapbuf_size5_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_46_sram;
wire [0:2] mux_tree_tapbuf_size5_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_47_sram;
wire [0:2] mux_tree_tapbuf_size5_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_48_sram;
wire [0:2] mux_tree_tapbuf_size5_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_49_sram;
wire [0:2] mux_tree_tapbuf_size5_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_50_sram;
wire [0:2] mux_tree_tapbuf_size5_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_51_sram;
wire [0:2] mux_tree_tapbuf_size5_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_52_sram;
wire [0:2] mux_tree_tapbuf_size5_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_53_sram;
wire [0:2] mux_tree_tapbuf_size5_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_54_sram;
wire [0:2] mux_tree_tapbuf_size5_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_55_sram;
wire [0:2] mux_tree_tapbuf_size5_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_56_sram;
wire [0:2] mux_tree_tapbuf_size5_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_57_sram;
wire [0:2] mux_tree_tapbuf_size5_57_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_58_sram;
wire [0:2] mux_tree_tapbuf_size5_58_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_59_sram;
wire [0:2] mux_tree_tapbuf_size5_59_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_60_sram;
wire [0:2] mux_tree_tapbuf_size5_60_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_61_sram;
wire [0:2] mux_tree_tapbuf_size5_61_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_62_sram;
wire [0:2] mux_tree_tapbuf_size5_62_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_63_sram;
wire [0:2] mux_tree_tapbuf_size5_63_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_64_sram;
wire [0:2] mux_tree_tapbuf_size5_64_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_65_sram;
wire [0:2] mux_tree_tapbuf_size5_65_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_66_sram;
wire [0:2] mux_tree_tapbuf_size5_66_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_67_sram;
wire [0:2] mux_tree_tapbuf_size5_67_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_68_sram;
wire [0:2] mux_tree_tapbuf_size5_68_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_69_sram;
wire [0:2] mux_tree_tapbuf_size5_69_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_70_sram;
wire [0:2] mux_tree_tapbuf_size5_70_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_71_sram;
wire [0:2] mux_tree_tapbuf_size5_71_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_72_sram;
wire [0:2] mux_tree_tapbuf_size5_72_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_73_sram;
wire [0:2] mux_tree_tapbuf_size5_73_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_74_sram;
wire [0:2] mux_tree_tapbuf_size5_74_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_75_sram;
wire [0:2] mux_tree_tapbuf_size5_75_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_76_sram;
wire [0:2] mux_tree_tapbuf_size5_76_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_77_sram;
wire [0:2] mux_tree_tapbuf_size5_77_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_78_sram;
wire [0:2] mux_tree_tapbuf_size5_78_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_79_sram;
wire [0:2] mux_tree_tapbuf_size5_79_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_80_sram;
wire [0:2] mux_tree_tapbuf_size5_80_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_11_sram;
wire [0:2] mux_tree_tapbuf_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_12_sram;
wire [0:2] mux_tree_tapbuf_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_13_sram;
wire [0:2] mux_tree_tapbuf_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_14_sram;
wire [0:2] mux_tree_tapbuf_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_15_sram;
wire [0:2] mux_tree_tapbuf_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_16_sram;
wire [0:2] mux_tree_tapbuf_size6_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_17_sram;
wire [0:2] mux_tree_tapbuf_size6_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_18_sram;
wire [0:2] mux_tree_tapbuf_size6_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_19_sram;
wire [0:2] mux_tree_tapbuf_size6_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_20_sram;
wire [0:2] mux_tree_tapbuf_size6_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_21_sram;
wire [0:2] mux_tree_tapbuf_size6_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_22_sram;
wire [0:2] mux_tree_tapbuf_size6_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_23_sram;
wire [0:2] mux_tree_tapbuf_size6_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_24_sram;
wire [0:2] mux_tree_tapbuf_size6_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_25_sram;
wire [0:2] mux_tree_tapbuf_size6_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_26_sram;
wire [0:2] mux_tree_tapbuf_size6_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_27_sram;
wire [0:2] mux_tree_tapbuf_size6_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_28_sram;
wire [0:2] mux_tree_tapbuf_size6_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_29_sram;
wire [0:2] mux_tree_tapbuf_size6_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_30_sram;
wire [0:2] mux_tree_tapbuf_size6_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_31_sram;
wire [0:2] mux_tree_tapbuf_size6_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_32_sram;
wire [0:2] mux_tree_tapbuf_size6_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_33_sram;
wire [0:2] mux_tree_tapbuf_size6_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_34_sram;
wire [0:2] mux_tree_tapbuf_size6_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_35_sram;
wire [0:2] mux_tree_tapbuf_size6_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_36_sram;
wire [0:2] mux_tree_tapbuf_size6_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_37_sram;
wire [0:2] mux_tree_tapbuf_size6_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_38_sram;
wire [0:2] mux_tree_tapbuf_size6_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_39_sram;
wire [0:2] mux_tree_tapbuf_size6_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_40_sram;
wire [0:2] mux_tree_tapbuf_size6_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_41_sram;
wire [0:2] mux_tree_tapbuf_size6_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_42_sram;
wire [0:2] mux_tree_tapbuf_size6_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_43_sram;
wire [0:2] mux_tree_tapbuf_size6_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_44_sram;
wire [0:2] mux_tree_tapbuf_size6_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_45_sram;
wire [0:2] mux_tree_tapbuf_size6_45_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_46_sram;
wire [0:2] mux_tree_tapbuf_size6_46_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_47_sram;
wire [0:2] mux_tree_tapbuf_size6_47_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_48_sram;
wire [0:2] mux_tree_tapbuf_size6_48_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_49_sram;
wire [0:2] mux_tree_tapbuf_size6_49_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_50_sram;
wire [0:2] mux_tree_tapbuf_size6_50_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_51_sram;
wire [0:2] mux_tree_tapbuf_size6_51_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_52_sram;
wire [0:2] mux_tree_tapbuf_size6_52_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_53_sram;
wire [0:2] mux_tree_tapbuf_size6_53_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_54_sram;
wire [0:2] mux_tree_tapbuf_size6_54_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_55_sram;
wire [0:2] mux_tree_tapbuf_size6_55_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_56_sram;
wire [0:2] mux_tree_tapbuf_size6_56_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_4_sram;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_5_sram;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_6_sram;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_7_sram;
wire [0:2] mux_tree_tapbuf_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_8_sram;
wire [0:2] mux_tree_tapbuf_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_9_sram;
wire [0:2] mux_tree_tapbuf_size7_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[193] = chany_top_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[194] = chany_top_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[195] = chany_top_in[194];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[197] = chany_top_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[198] = chany_top_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[199] = chany_top_in[198];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[201] = chany_top_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[202] = chany_top_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[203] = chany_top_in[202];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[205] = chany_top_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[206] = chany_top_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[207] = chany_top_in[206];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[209] = chany_top_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[210] = chany_top_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[211] = chany_top_in[210];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[213] = chany_top_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[214] = chany_top_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[215] = chany_top_in[214];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[217] = chany_top_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[218] = chany_top_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[219] = chany_top_in[218];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[221] = chany_top_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[222] = chany_top_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[223] = chany_top_in[222];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[225] = chany_top_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[226] = chany_top_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[227] = chany_top_in[226];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[229] = chany_top_in[228];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[230] = chany_top_in[229];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[231] = chany_top_in[230];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[233] = chany_top_in[232];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[234] = chany_top_in[233];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[235] = chany_top_in[234];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[237] = chany_top_in[236];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[238] = chany_top_in[237];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[239] = chany_top_in[238];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[241] = chany_top_in[240];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[242] = chany_top_in[241];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[243] = chany_top_in[242];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[245] = chany_top_in[244];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[246] = chany_top_in[245];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[247] = chany_top_in[246];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[249] = chany_top_in[248];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[250] = chany_top_in[249];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[251] = chany_top_in[250];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[253] = chany_top_in[252];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[254] = chany_top_in[253];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[255] = chany_top_in[254];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[257] = chany_top_in[256];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[258] = chany_top_in[257];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[259] = chany_top_in[258];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[261] = chany_top_in[260];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[262] = chany_top_in[261];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[263] = chany_top_in[262];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[265] = chany_top_in[264];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[266] = chany_top_in[265];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[267] = chany_top_in[266];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[269] = chany_top_in[268];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[270] = chany_top_in[269];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[271] = chany_top_in[270];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[273] = chany_top_in[272];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[274] = chany_top_in[273];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[275] = chany_top_in[274];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[277] = chany_top_in[276];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[278] = chany_top_in[277];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[279] = chany_top_in[278];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[281] = chany_top_in[280];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[282] = chany_top_in[281];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[283] = chany_top_in[282];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[285] = chany_top_in[284];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[286] = chany_top_in[285];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[287] = chany_top_in[286];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[289] = chany_top_in[288];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[290] = chany_top_in[289];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[291] = chany_top_in[290];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[293] = chany_top_in[292];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[294] = chany_top_in[293];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[295] = chany_top_in[294];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 32 -----
	assign chanx_right_out[295] = right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_[0];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 611 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 615 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 619 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 623 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 627 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 631 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 635 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 639 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 643 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 647 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 651 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 655 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 659 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 663 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 667 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 671 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 675 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 679 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 683 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 687 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 691 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 695 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 699 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 703 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 707 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 711 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 714 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 715 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 718 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 719 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 722 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 723 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 726 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 727 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 730 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 731 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 734 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 735 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 738 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 739 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 742 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 743 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 746 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 747 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 750 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 751 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 754 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 755 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 758 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 759 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 762 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 763 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 766 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 767 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 770 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 771 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 774 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 775 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 778 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 779 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 782 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 783 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 786 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 787 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 791 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 792 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 795 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 796 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 799 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 800 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[193] = chany_bottom_in[192];
// ----- Local connection due to Wire 803 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[194] = chany_bottom_in[193];
// ----- Local connection due to Wire 804 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[195] = chany_bottom_in[194];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chany_bottom_in[196];
// ----- Local connection due to Wire 807 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[198] = chany_bottom_in[197];
// ----- Local connection due to Wire 808 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[199] = chany_bottom_in[198];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[201] = chany_bottom_in[200];
// ----- Local connection due to Wire 811 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[202] = chany_bottom_in[201];
// ----- Local connection due to Wire 812 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[203] = chany_bottom_in[202];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[205] = chany_bottom_in[204];
// ----- Local connection due to Wire 815 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chany_bottom_in[205];
// ----- Local connection due to Wire 816 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[207] = chany_bottom_in[206];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[209] = chany_bottom_in[208];
// ----- Local connection due to Wire 819 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[210] = chany_bottom_in[209];
// ----- Local connection due to Wire 820 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[211] = chany_bottom_in[210];
// ----- Local connection due to Wire 822 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[213] = chany_bottom_in[212];
// ----- Local connection due to Wire 823 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[214] = chany_bottom_in[213];
// ----- Local connection due to Wire 824 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chany_bottom_in[214];
// ----- Local connection due to Wire 826 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[217] = chany_bottom_in[216];
// ----- Local connection due to Wire 827 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[218] = chany_bottom_in[217];
// ----- Local connection due to Wire 828 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[219] = chany_bottom_in[218];
// ----- Local connection due to Wire 830 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[221] = chany_bottom_in[220];
// ----- Local connection due to Wire 831 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[222] = chany_bottom_in[221];
// ----- Local connection due to Wire 832 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[223] = chany_bottom_in[222];
// ----- Local connection due to Wire 834 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[225] = chany_bottom_in[224];
// ----- Local connection due to Wire 835 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[226] = chany_bottom_in[225];
// ----- Local connection due to Wire 836 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[227] = chany_bottom_in[226];
// ----- Local connection due to Wire 838 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[229] = chany_bottom_in[228];
// ----- Local connection due to Wire 839 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[230] = chany_bottom_in[229];
// ----- Local connection due to Wire 840 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[231] = chany_bottom_in[230];
// ----- Local connection due to Wire 842 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[233] = chany_bottom_in[232];
// ----- Local connection due to Wire 843 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[234] = chany_bottom_in[233];
// ----- Local connection due to Wire 844 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[235] = chany_bottom_in[234];
// ----- Local connection due to Wire 846 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[237] = chany_bottom_in[236];
// ----- Local connection due to Wire 847 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[238] = chany_bottom_in[237];
// ----- Local connection due to Wire 848 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[239] = chany_bottom_in[238];
// ----- Local connection due to Wire 850 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[241] = chany_bottom_in[240];
// ----- Local connection due to Wire 851 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[242] = chany_bottom_in[241];
// ----- Local connection due to Wire 852 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[243] = chany_bottom_in[242];
// ----- Local connection due to Wire 854 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[245] = chany_bottom_in[244];
// ----- Local connection due to Wire 855 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[246] = chany_bottom_in[245];
// ----- Local connection due to Wire 856 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[247] = chany_bottom_in[246];
// ----- Local connection due to Wire 858 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[249] = chany_bottom_in[248];
// ----- Local connection due to Wire 859 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[250] = chany_bottom_in[249];
// ----- Local connection due to Wire 860 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[251] = chany_bottom_in[250];
// ----- Local connection due to Wire 862 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[253] = chany_bottom_in[252];
// ----- Local connection due to Wire 863 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[254] = chany_bottom_in[253];
// ----- Local connection due to Wire 864 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[255] = chany_bottom_in[254];
// ----- Local connection due to Wire 866 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[257] = chany_bottom_in[256];
// ----- Local connection due to Wire 867 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[258] = chany_bottom_in[257];
// ----- Local connection due to Wire 868 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[259] = chany_bottom_in[258];
// ----- Local connection due to Wire 870 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[261] = chany_bottom_in[260];
// ----- Local connection due to Wire 871 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[262] = chany_bottom_in[261];
// ----- Local connection due to Wire 872 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[263] = chany_bottom_in[262];
// ----- Local connection due to Wire 874 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[265] = chany_bottom_in[264];
// ----- Local connection due to Wire 875 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[266] = chany_bottom_in[265];
// ----- Local connection due to Wire 876 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[267] = chany_bottom_in[266];
// ----- Local connection due to Wire 878 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[269] = chany_bottom_in[268];
// ----- Local connection due to Wire 879 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[270] = chany_bottom_in[269];
// ----- Local connection due to Wire 880 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[271] = chany_bottom_in[270];
// ----- Local connection due to Wire 882 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[273] = chany_bottom_in[272];
// ----- Local connection due to Wire 883 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[274] = chany_bottom_in[273];
// ----- Local connection due to Wire 884 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[275] = chany_bottom_in[274];
// ----- Local connection due to Wire 886 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[277] = chany_bottom_in[276];
// ----- Local connection due to Wire 887 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[278] = chany_bottom_in[277];
// ----- Local connection due to Wire 888 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[279] = chany_bottom_in[278];
// ----- Local connection due to Wire 890 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[281] = chany_bottom_in[280];
// ----- Local connection due to Wire 891 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[282] = chany_bottom_in[281];
// ----- Local connection due to Wire 892 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[283] = chany_bottom_in[282];
// ----- Local connection due to Wire 894 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[285] = chany_bottom_in[284];
// ----- Local connection due to Wire 895 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[286] = chany_bottom_in[285];
// ----- Local connection due to Wire 896 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[287] = chany_bottom_in[286];
// ----- Local connection due to Wire 898 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[289] = chany_bottom_in[288];
// ----- Local connection due to Wire 899 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[290] = chany_bottom_in[289];
// ----- Local connection due to Wire 900 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[291] = chany_bottom_in[290];
// ----- Local connection due to Wire 902 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[293] = chany_bottom_in[292];
// ----- Local connection due to Wire 903 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[294] = chany_bottom_in[293];
// ----- Local connection due to Wire 904 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[295] = chany_bottom_in[294];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size6 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[1], chanx_right_in[75], chanx_right_in[149], chanx_right_in[223]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size6 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[2], chanx_right_in[76], chanx_right_in[150], chanx_right_in[224]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size6 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[3], chanx_right_in[77], chanx_right_in[151], chanx_right_in[225]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size6 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[4], chanx_right_in[78], chanx_right_in[152], chanx_right_in[226]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size6 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[5], chanx_right_in[79], chanx_right_in[153], chanx_right_in[227]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size6 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[6], chanx_right_in[80], chanx_right_in[154], chanx_right_in[228]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size6 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[7], chanx_right_in[81], chanx_right_in[155], chanx_right_in[229]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_41 (
		.in({chanx_right_in[67], chanx_right_in[141], chanx_right_in[215], chanx_right_in[289], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size6 mux_bottom_track_49 (
		.in({chanx_right_in[66], chanx_right_in[140], chanx_right_in[214], chanx_right_in[288], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_57 (
		.in({chanx_right_in[65], chanx_right_in[139], chanx_right_in[213], chanx_right_in[287], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size6 mux_bottom_track_65 (
		.in({chanx_right_in[64], chanx_right_in[138], chanx_right_in[212], chanx_right_in[286], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size6 mux_bottom_track_113 (
		.in({chanx_right_in[58], chanx_right_in[132], chanx_right_in[206], chanx_right_in[280], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_11_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size6 mux_bottom_track_121 (
		.in({chanx_right_in[57], chanx_right_in[131], chanx_right_in[205], chanx_right_in[279], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_12_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size6 mux_bottom_track_145 (
		.in({chanx_right_in[54], chanx_right_in[128], chanx_right_in[202], chanx_right_in[276], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_13_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size6 mux_bottom_track_153 (
		.in({chanx_right_in[53], chanx_right_in[127], chanx_right_in[201], chanx_right_in[275], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_14_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size6 mux_bottom_track_161 (
		.in({chanx_right_in[52], chanx_right_in[126], chanx_right_in[200], chanx_right_in[274], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_15_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size6 mux_bottom_track_169 (
		.in({chanx_right_in[51], chanx_right_in[125], chanx_right_in[199], chanx_right_in[273], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_16_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size6 mux_bottom_track_177 (
		.in({chanx_right_in[50], chanx_right_in[124], chanx_right_in[198], chanx_right_in[272], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_17_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size6 mux_bottom_track_185 (
		.in({chanx_right_in[49], chanx_right_in[123], chanx_right_in[197], chanx_right_in[271], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_18_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size6 mux_bottom_track_193 (
		.in({chanx_right_in[48], chanx_right_in[122], chanx_right_in[196], chanx_right_in[270], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_19_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size6 mux_bottom_track_217 (
		.in({chanx_right_in[45], chanx_right_in[119], chanx_right_in[193], chanx_right_in[267], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_20_sram_inv[0:2]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size6 mux_bottom_track_225 (
		.in({chanx_right_in[44], chanx_right_in[118], chanx_right_in[192], chanx_right_in[266], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_21_sram_inv[0:2]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size6 mux_bottom_track_233 (
		.in({chanx_right_in[43], chanx_right_in[117], chanx_right_in[191], chanx_right_in[265], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_22_sram_inv[0:2]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size6 mux_bottom_track_241 (
		.in({chanx_right_in[42], chanx_right_in[116], chanx_right_in[190], chanx_right_in[264], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_23_sram_inv[0:2]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size6 mux_bottom_track_249 (
		.in({chanx_right_in[41], chanx_right_in[115], chanx_right_in[189], chanx_right_in[263], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_24_sram_inv[0:2]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size6 mux_bottom_track_257 (
		.in({chanx_right_in[40], chanx_right_in[114], chanx_right_in[188], chanx_right_in[262], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_25_sram_inv[0:2]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size6 mux_bottom_track_265 (
		.in({chanx_right_in[39], chanx_right_in[113], chanx_right_in[187], chanx_right_in[261], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_26_sram_inv[0:2]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size6 mux_bottom_track_289 (
		.in({chanx_right_in[36], chanx_right_in[110], chanx_right_in[184], chanx_right_in[258], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_27_sram_inv[0:2]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size6 mux_bottom_track_297 (
		.in({chanx_right_in[35], chanx_right_in[109], chanx_right_in[183], chanx_right_in[257], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_28_sram_inv[0:2]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size6 mux_bottom_track_305 (
		.in({chanx_right_in[34], chanx_right_in[108], chanx_right_in[182], chanx_right_in[256], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_29_sram_inv[0:2]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size6 mux_bottom_track_313 (
		.in({chanx_right_in[33], chanx_right_in[107], chanx_right_in[181], chanx_right_in[255], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_30_sram_inv[0:2]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size6 mux_bottom_track_321 (
		.in({chanx_right_in[32], chanx_right_in[106], chanx_right_in[180], chanx_right_in[254], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_31_sram_inv[0:2]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size6 mux_bottom_track_329 (
		.in({chanx_right_in[31], chanx_right_in[105], chanx_right_in[179], chanx_right_in[253], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_32_sram_inv[0:2]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size6 mux_bottom_track_337 (
		.in({chanx_right_in[30], chanx_right_in[104], chanx_right_in[178], chanx_right_in[252], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_33_sram_inv[0:2]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size6 mux_bottom_track_361 (
		.in({chanx_right_in[27], chanx_right_in[101], chanx_right_in[175], chanx_right_in[249], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_34_sram_inv[0:2]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size6 mux_bottom_track_369 (
		.in({chanx_right_in[26], chanx_right_in[100], chanx_right_in[174], chanx_right_in[248], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_35_sram_inv[0:2]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size6 mux_bottom_track_377 (
		.in({chanx_right_in[25], chanx_right_in[99], chanx_right_in[173], chanx_right_in[247], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_36_sram_inv[0:2]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size6 mux_bottom_track_385 (
		.in({chanx_right_in[24], chanx_right_in[98], chanx_right_in[172], chanx_right_in[246], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_37_sram_inv[0:2]),
		.out(chany_bottom_out[192]));

	mux_tree_tapbuf_size6 mux_bottom_track_393 (
		.in({chanx_right_in[23], chanx_right_in[97], chanx_right_in[171], chanx_right_in[245], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_38_sram_inv[0:2]),
		.out(chany_bottom_out[196]));

	mux_tree_tapbuf_size6 mux_bottom_track_401 (
		.in({chanx_right_in[22], chanx_right_in[96], chanx_right_in[170], chanx_right_in[244], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_39_sram_inv[0:2]),
		.out(chany_bottom_out[200]));

	mux_tree_tapbuf_size6 mux_bottom_track_409 (
		.in({chanx_right_in[21], chanx_right_in[95], chanx_right_in[169], chanx_right_in[243], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_40_sram_inv[0:2]),
		.out(chany_bottom_out[204]));

	mux_tree_tapbuf_size6 mux_bottom_track_433 (
		.in({chanx_right_in[18], chanx_right_in[92], chanx_right_in[166], chanx_right_in[240], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_41_sram_inv[0:2]),
		.out(chany_bottom_out[216]));

	mux_tree_tapbuf_size6 mux_bottom_track_441 (
		.in({chanx_right_in[17], chanx_right_in[91], chanx_right_in[165], chanx_right_in[239], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_42_sram_inv[0:2]),
		.out(chany_bottom_out[220]));

	mux_tree_tapbuf_size6 mux_bottom_track_449 (
		.in({chanx_right_in[16], chanx_right_in[90], chanx_right_in[164], chanx_right_in[238], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_43_sram_inv[0:2]),
		.out(chany_bottom_out[224]));

	mux_tree_tapbuf_size6 mux_bottom_track_457 (
		.in({chanx_right_in[15], chanx_right_in[89], chanx_right_in[163], chanx_right_in[237], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_44_sram_inv[0:2]),
		.out(chany_bottom_out[228]));

	mux_tree_tapbuf_size6 mux_bottom_track_465 (
		.in({chanx_right_in[14], chanx_right_in[88], chanx_right_in[162], chanx_right_in[236], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_45_sram_inv[0:2]),
		.out(chany_bottom_out[232]));

	mux_tree_tapbuf_size6 mux_bottom_track_473 (
		.in({chanx_right_in[13], chanx_right_in[87], chanx_right_in[161], chanx_right_in[235], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_46_sram_inv[0:2]),
		.out(chany_bottom_out[236]));

	mux_tree_tapbuf_size6 mux_bottom_track_481 (
		.in({chanx_right_in[12], chanx_right_in[86], chanx_right_in[160], chanx_right_in[234], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_47_sram_inv[0:2]),
		.out(chany_bottom_out[240]));

	mux_tree_tapbuf_size6 mux_bottom_track_505 (
		.in({chanx_right_in[9], chanx_right_in[83], chanx_right_in[157], chanx_right_in[231], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_48_sram_inv[0:2]),
		.out(chany_bottom_out[252]));

	mux_tree_tapbuf_size6 mux_bottom_track_513 (
		.in({chanx_right_in[8], chanx_right_in[82], chanx_right_in[156], chanx_right_in[230], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_49_sram_inv[0:2]),
		.out(chany_bottom_out[256]));

	mux_tree_tapbuf_size6 mux_bottom_track_521 (
		.in({chanx_right_in[7], chanx_right_in[81], chanx_right_in[155], chanx_right_in[229], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_50_sram_inv[0:2]),
		.out(chany_bottom_out[260]));

	mux_tree_tapbuf_size6 mux_bottom_track_529 (
		.in({chanx_right_in[6], chanx_right_in[80], chanx_right_in[154], chanx_right_in[228], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_51_sram_inv[0:2]),
		.out(chany_bottom_out[264]));

	mux_tree_tapbuf_size6 mux_bottom_track_537 (
		.in({chanx_right_in[5], chanx_right_in[79], chanx_right_in[153], chanx_right_in[227], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_52_sram_inv[0:2]),
		.out(chany_bottom_out[268]));

	mux_tree_tapbuf_size6 mux_bottom_track_545 (
		.in({chanx_right_in[4], chanx_right_in[78], chanx_right_in[152], chanx_right_in[226], bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_53_sram_inv[0:2]),
		.out(chany_bottom_out[272]));

	mux_tree_tapbuf_size6 mux_bottom_track_553 (
		.in({chanx_right_in[3], chanx_right_in[77], chanx_right_in[151], chanx_right_in[225], bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_54_sram_inv[0:2]),
		.out(chany_bottom_out[276]));

	mux_tree_tapbuf_size6 mux_bottom_track_577 (
		.in({chanx_right_in[0], chanx_right_in[74], chanx_right_in[148], chanx_right_in[222], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_55_sram_inv[0:2]),
		.out(chany_bottom_out[288]));

	mux_tree_tapbuf_size6 mux_bottom_track_585 (
		.in({chanx_right_in[73], chanx_right_in[147], chanx_right_in[221], chanx_right_in[295], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_56_sram_inv[0:2]),
		.out(chany_bottom_out[292]));

	mux_tree_tapbuf_size6_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_16_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_17_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_18_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_19_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_20_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_21_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_22_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_23_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_24_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_25_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_26_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_27_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_28_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_29_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_30_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_31_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_32_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_33_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_34_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_35_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_36_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_37_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_38_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_39_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_40_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_41_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_42_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_43_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_44_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_45_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_46_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_47_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_48_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_49_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_50_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_51_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_52_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_53_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_54_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_577 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_55_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_585 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_55_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_56_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[8], chanx_right_in[82], chanx_right_in[156], chanx_right_in[230]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size5 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[9], chanx_right_in[83], chanx_right_in[157], chanx_right_in[231]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size5 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[10], chanx_right_in[84], chanx_right_in[158], chanx_right_in[232]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size5 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[11], chanx_right_in[85], chanx_right_in[159], chanx_right_in[233]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size5 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[12], chanx_right_in[86], chanx_right_in[160], chanx_right_in[234]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size5 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[13], chanx_right_in[87], chanx_right_in[161], chanx_right_in[235]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size5 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[14], chanx_right_in[88], chanx_right_in[162], chanx_right_in[236]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size5 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[15], chanx_right_in[89], chanx_right_in[163], chanx_right_in[237]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size5 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[16], chanx_right_in[90], chanx_right_in[164], chanx_right_in[238]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size5 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[17], chanx_right_in[91], chanx_right_in[165], chanx_right_in[239]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size5 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[18], chanx_right_in[92], chanx_right_in[166], chanx_right_in[240]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size5 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[19], chanx_right_in[93], chanx_right_in[167], chanx_right_in[241]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size5 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[20], chanx_right_in[94], chanx_right_in[168], chanx_right_in[242]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size5 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[21], chanx_right_in[95], chanx_right_in[169], chanx_right_in[243]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size5 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[22], chanx_right_in[96], chanx_right_in[170], chanx_right_in[244]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size5 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[23], chanx_right_in[97], chanx_right_in[171], chanx_right_in[245]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size5 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[24], chanx_right_in[98], chanx_right_in[172], chanx_right_in[246]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size5 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[25], chanx_right_in[99], chanx_right_in[173], chanx_right_in[247]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size5 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[26], chanx_right_in[100], chanx_right_in[174], chanx_right_in[248]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size5 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[27], chanx_right_in[101], chanx_right_in[175], chanx_right_in[249]}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size5 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[28], chanx_right_in[102], chanx_right_in[176], chanx_right_in[250]}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size5 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[29], chanx_right_in[103], chanx_right_in[177], chanx_right_in[251]}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size5 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[30], chanx_right_in[104], chanx_right_in[178], chanx_right_in[252]}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size5 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[31], chanx_right_in[105], chanx_right_in[179], chanx_right_in[253]}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size5 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[32], chanx_right_in[106], chanx_right_in[180], chanx_right_in[254]}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size5 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[33], chanx_right_in[107], chanx_right_in[181], chanx_right_in[255]}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size5 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[34], chanx_right_in[108], chanx_right_in[182], chanx_right_in[256]}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size5 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[35], chanx_right_in[109], chanx_right_in[183], chanx_right_in[257]}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size5 mux_top_track_280 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[36], chanx_right_in[110], chanx_right_in[184], chanx_right_in[258]}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size5 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[37], chanx_right_in[111], chanx_right_in[185], chanx_right_in[259]}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size5 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[38], chanx_right_in[112], chanx_right_in[186], chanx_right_in[260]}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size5 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[39], chanx_right_in[113], chanx_right_in[187], chanx_right_in[261]}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size5 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[40], chanx_right_in[114], chanx_right_in[188], chanx_right_in[262]}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size5 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[41], chanx_right_in[115], chanx_right_in[189], chanx_right_in[263]}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size5 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[42], chanx_right_in[116], chanx_right_in[190], chanx_right_in[264]}),
		.sram(mux_tree_tapbuf_size5_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_34_sram_inv[0:2]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size5 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[43], chanx_right_in[117], chanx_right_in[191], chanx_right_in[265]}),
		.sram(mux_tree_tapbuf_size5_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_35_sram_inv[0:2]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size5 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[44], chanx_right_in[118], chanx_right_in[192], chanx_right_in[266]}),
		.sram(mux_tree_tapbuf_size5_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_36_sram_inv[0:2]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size5 mux_top_track_352 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[45], chanx_right_in[119], chanx_right_in[193], chanx_right_in[267]}),
		.sram(mux_tree_tapbuf_size5_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_37_sram_inv[0:2]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size5 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[46], chanx_right_in[120], chanx_right_in[194], chanx_right_in[268]}),
		.sram(mux_tree_tapbuf_size5_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_38_sram_inv[0:2]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size5 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[47], chanx_right_in[121], chanx_right_in[195], chanx_right_in[269]}),
		.sram(mux_tree_tapbuf_size5_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_39_sram_inv[0:2]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size5 mux_top_track_376 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[48], chanx_right_in[122], chanx_right_in[196], chanx_right_in[270]}),
		.sram(mux_tree_tapbuf_size5_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_40_sram_inv[0:2]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size5 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[49], chanx_right_in[123], chanx_right_in[197], chanx_right_in[271]}),
		.sram(mux_tree_tapbuf_size5_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_41_sram_inv[0:2]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size5 mux_top_track_392 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[50], chanx_right_in[124], chanx_right_in[198], chanx_right_in[272]}),
		.sram(mux_tree_tapbuf_size5_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_42_sram_inv[0:2]),
		.out(chany_top_out[196]));

	mux_tree_tapbuf_size5 mux_top_track_400 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[51], chanx_right_in[125], chanx_right_in[199], chanx_right_in[273]}),
		.sram(mux_tree_tapbuf_size5_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_43_sram_inv[0:2]),
		.out(chany_top_out[200]));

	mux_tree_tapbuf_size5 mux_top_track_408 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[52], chanx_right_in[126], chanx_right_in[200], chanx_right_in[274]}),
		.sram(mux_tree_tapbuf_size5_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_44_sram_inv[0:2]),
		.out(chany_top_out[204]));

	mux_tree_tapbuf_size5 mux_top_track_416 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[53], chanx_right_in[127], chanx_right_in[201], chanx_right_in[275]}),
		.sram(mux_tree_tapbuf_size5_45_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_45_sram_inv[0:2]),
		.out(chany_top_out[208]));

	mux_tree_tapbuf_size5 mux_top_track_424 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[54], chanx_right_in[128], chanx_right_in[202], chanx_right_in[276]}),
		.sram(mux_tree_tapbuf_size5_46_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_46_sram_inv[0:2]),
		.out(chany_top_out[212]));

	mux_tree_tapbuf_size5 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[55], chanx_right_in[129], chanx_right_in[203], chanx_right_in[277]}),
		.sram(mux_tree_tapbuf_size5_47_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_47_sram_inv[0:2]),
		.out(chany_top_out[216]));

	mux_tree_tapbuf_size5 mux_top_track_440 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[56], chanx_right_in[130], chanx_right_in[204], chanx_right_in[278]}),
		.sram(mux_tree_tapbuf_size5_48_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_48_sram_inv[0:2]),
		.out(chany_top_out[220]));

	mux_tree_tapbuf_size5 mux_top_track_448 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[57], chanx_right_in[131], chanx_right_in[205], chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size5_49_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_49_sram_inv[0:2]),
		.out(chany_top_out[224]));

	mux_tree_tapbuf_size5 mux_top_track_456 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[58], chanx_right_in[132], chanx_right_in[206], chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size5_50_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_50_sram_inv[0:2]),
		.out(chany_top_out[228]));

	mux_tree_tapbuf_size5 mux_top_track_464 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[59], chanx_right_in[133], chanx_right_in[207], chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size5_51_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_51_sram_inv[0:2]),
		.out(chany_top_out[232]));

	mux_tree_tapbuf_size5 mux_top_track_472 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[60], chanx_right_in[134], chanx_right_in[208], chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size5_52_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_52_sram_inv[0:2]),
		.out(chany_top_out[236]));

	mux_tree_tapbuf_size5 mux_top_track_480 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[61], chanx_right_in[135], chanx_right_in[209], chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size5_53_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_53_sram_inv[0:2]),
		.out(chany_top_out[240]));

	mux_tree_tapbuf_size5 mux_top_track_488 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[62], chanx_right_in[136], chanx_right_in[210], chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size5_54_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_54_sram_inv[0:2]),
		.out(chany_top_out[244]));

	mux_tree_tapbuf_size5 mux_top_track_496 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[63], chanx_right_in[137], chanx_right_in[211], chanx_right_in[285]}),
		.sram(mux_tree_tapbuf_size5_55_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_55_sram_inv[0:2]),
		.out(chany_top_out[248]));

	mux_tree_tapbuf_size5 mux_top_track_504 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[64], chanx_right_in[138], chanx_right_in[212], chanx_right_in[286]}),
		.sram(mux_tree_tapbuf_size5_56_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_56_sram_inv[0:2]),
		.out(chany_top_out[252]));

	mux_tree_tapbuf_size5 mux_top_track_512 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[65], chanx_right_in[139], chanx_right_in[213], chanx_right_in[287]}),
		.sram(mux_tree_tapbuf_size5_57_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_57_sram_inv[0:2]),
		.out(chany_top_out[256]));

	mux_tree_tapbuf_size5 mux_top_track_520 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[66], chanx_right_in[140], chanx_right_in[214], chanx_right_in[288]}),
		.sram(mux_tree_tapbuf_size5_58_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_58_sram_inv[0:2]),
		.out(chany_top_out[260]));

	mux_tree_tapbuf_size5 mux_top_track_528 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[67], chanx_right_in[141], chanx_right_in[215], chanx_right_in[289]}),
		.sram(mux_tree_tapbuf_size5_59_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_59_sram_inv[0:2]),
		.out(chany_top_out[264]));

	mux_tree_tapbuf_size5 mux_top_track_536 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[68], chanx_right_in[142], chanx_right_in[216], chanx_right_in[290]}),
		.sram(mux_tree_tapbuf_size5_60_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_60_sram_inv[0:2]),
		.out(chany_top_out[268]));

	mux_tree_tapbuf_size5 mux_top_track_544 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[69], chanx_right_in[143], chanx_right_in[217], chanx_right_in[291]}),
		.sram(mux_tree_tapbuf_size5_61_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_61_sram_inv[0:2]),
		.out(chany_top_out[272]));

	mux_tree_tapbuf_size5 mux_top_track_552 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[70], chanx_right_in[144], chanx_right_in[218], chanx_right_in[292]}),
		.sram(mux_tree_tapbuf_size5_62_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_62_sram_inv[0:2]),
		.out(chany_top_out[276]));

	mux_tree_tapbuf_size5 mux_top_track_560 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[71], chanx_right_in[145], chanx_right_in[219], chanx_right_in[293]}),
		.sram(mux_tree_tapbuf_size5_63_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_63_sram_inv[0:2]),
		.out(chany_top_out[280]));

	mux_tree_tapbuf_size5 mux_top_track_568 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[72], chanx_right_in[146], chanx_right_in[220], chanx_right_in[294]}),
		.sram(mux_tree_tapbuf_size5_64_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_64_sram_inv[0:2]),
		.out(chany_top_out[284]));

	mux_tree_tapbuf_size5 mux_top_track_576 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[73], chanx_right_in[147], chanx_right_in[221], chanx_right_in[295]}),
		.sram(mux_tree_tapbuf_size5_65_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_65_sram_inv[0:2]),
		.out(chany_top_out[288]));

	mux_tree_tapbuf_size5 mux_top_track_584 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[0], chanx_right_in[74], chanx_right_in[148], chanx_right_in[222]}),
		.sram(mux_tree_tapbuf_size5_66_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_66_sram_inv[0:2]),
		.out(chany_top_out[292]));

	mux_tree_tapbuf_size5 mux_bottom_track_129 (
		.in({chanx_right_in[56], chanx_right_in[130], chanx_right_in[204], chanx_right_in[278], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_67_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_67_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size5 mux_bottom_track_137 (
		.in({chanx_right_in[55], chanx_right_in[129], chanx_right_in[203], chanx_right_in[277], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_68_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_68_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size5 mux_bottom_track_201 (
		.in({chanx_right_in[47], chanx_right_in[121], chanx_right_in[195], chanx_right_in[269], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_69_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_69_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size5 mux_bottom_track_209 (
		.in({chanx_right_in[46], chanx_right_in[120], chanx_right_in[194], chanx_right_in[268], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_70_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_70_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size5 mux_bottom_track_273 (
		.in({chanx_right_in[38], chanx_right_in[112], chanx_right_in[186], chanx_right_in[260], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_71_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_71_sram_inv[0:2]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size5 mux_bottom_track_281 (
		.in({chanx_right_in[37], chanx_right_in[111], chanx_right_in[185], chanx_right_in[259], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_72_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_72_sram_inv[0:2]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size5 mux_bottom_track_345 (
		.in({chanx_right_in[29], chanx_right_in[103], chanx_right_in[177], chanx_right_in[251], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_73_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_73_sram_inv[0:2]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size5 mux_bottom_track_353 (
		.in({chanx_right_in[28], chanx_right_in[102], chanx_right_in[176], chanx_right_in[250], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_74_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_74_sram_inv[0:2]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size5 mux_bottom_track_417 (
		.in({chanx_right_in[20], chanx_right_in[94], chanx_right_in[168], chanx_right_in[242], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_75_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_75_sram_inv[0:2]),
		.out(chany_bottom_out[208]));

	mux_tree_tapbuf_size5 mux_bottom_track_425 (
		.in({chanx_right_in[19], chanx_right_in[93], chanx_right_in[167], chanx_right_in[241], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_76_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_76_sram_inv[0:2]),
		.out(chany_bottom_out[212]));

	mux_tree_tapbuf_size5 mux_bottom_track_489 (
		.in({chanx_right_in[11], chanx_right_in[85], chanx_right_in[159], chanx_right_in[233], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_77_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_77_sram_inv[0:2]),
		.out(chany_bottom_out[244]));

	mux_tree_tapbuf_size5 mux_bottom_track_497 (
		.in({chanx_right_in[10], chanx_right_in[84], chanx_right_in[158], chanx_right_in[232], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_78_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_78_sram_inv[0:2]),
		.out(chany_bottom_out[248]));

	mux_tree_tapbuf_size5 mux_bottom_track_561 (
		.in({chanx_right_in[2], chanx_right_in[76], chanx_right_in[150], chanx_right_in[224], bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_79_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_79_sram_inv[0:2]),
		.out(chany_bottom_out[280]));

	mux_tree_tapbuf_size5 mux_bottom_track_569 (
		.in({chanx_right_in[1], chanx_right_in[75], chanx_right_in[149], chanx_right_in[223], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_80_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_80_sram_inv[0:2]),
		.out(chany_bottom_out[284]));

	mux_tree_tapbuf_size5_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_34_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_35_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_36_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_37_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_38_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_39_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_40_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_41_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_42_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_43_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_44_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_45_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_45_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_46_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_46_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_47_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_47_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_48_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_48_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_49_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_49_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_50_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_50_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_51_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_51_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_52_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_52_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_53_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_53_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_54_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_54_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_55_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_55_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_56_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_56_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_57_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_57_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_58_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_58_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_59_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_59_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_60_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_60_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_61_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_61_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_62_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_62_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_63_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_63_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_64_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_64_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_576 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_65_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_65_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_584 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_66_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_66_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_67_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_67_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_68_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_68_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_69_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_69_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_70_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_70_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_71_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_71_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_72_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_72_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_73_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_73_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_74_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_74_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_75_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_75_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_76_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_76_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_77_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_77_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_78_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_78_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_79_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_79_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_80_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_80_sram_inv[0:2]));

	mux_tree_tapbuf_size2 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size2_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size3 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size3 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size3 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size3 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size3 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size3 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size3 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size3 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size3 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size3 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size3 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size3 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size3 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size3 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size3 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size3 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[75], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size3 mux_right_track_40 (
		.in({chany_top_in[25], chany_top_in[79], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size3 mux_right_track_42 (
		.in({chany_top_in[26], chany_top_in[83], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size3 mux_right_track_44 (
		.in({chany_top_in[28], chany_top_in[87], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size3 mux_right_track_46 (
		.in({chany_top_in[29], chany_top_in[91], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size3 mux_right_track_48 (
		.in({chany_top_in[30], chany_top_in[95], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size3 mux_right_track_50 (
		.in({chany_top_in[32], chany_top_in[99], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size3 mux_right_track_52 (
		.in({chany_top_in[33], chany_top_in[103], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size3 mux_right_track_54 (
		.in({chany_top_in[34], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size3 mux_right_track_56 (
		.in({chany_top_in[36], chany_top_in[111], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size3 mux_right_track_58 (
		.in({chany_top_in[37], chany_top_in[115], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size3 mux_right_track_60 (
		.in({chany_top_in[38], chany_top_in[119], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size3 mux_right_track_62 (
		.in({chany_top_in[40], chany_top_in[123], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size3 mux_right_track_64 (
		.in({chany_top_in[41], chany_top_in[127], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size3 mux_right_track_66 (
		.in({chany_top_in[42], chany_top_in[131], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size3 mux_right_track_68 (
		.in({chany_top_in[44], chany_top_in[135], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size3 mux_right_track_70 (
		.in({chany_top_in[45], chany_top_in[139], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size3 mux_right_track_72 (
		.in({chany_top_in[46], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size3 mux_right_track_74 (
		.in({chany_top_in[48], chany_top_in[147], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size3 mux_right_track_76 (
		.in({chany_top_in[49], chany_top_in[151], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size3 mux_right_track_78 (
		.in({chany_top_in[50], chany_top_in[155], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size3 mux_right_track_80 (
		.in({chany_top_in[52], chany_top_in[159], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size3 mux_right_track_82 (
		.in({chany_top_in[53], chany_top_in[163], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size3 mux_right_track_84 (
		.in({chany_top_in[54], chany_top_in[167], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size3 mux_right_track_86 (
		.in({chany_top_in[56], chany_top_in[171], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size3 mux_right_track_88 (
		.in({chany_top_in[57], chany_top_in[175], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size3 mux_right_track_90 (
		.in({chany_top_in[58], chany_top_in[179], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size3 mux_right_track_92 (
		.in({chany_top_in[60], chany_top_in[183], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size3 mux_right_track_94 (
		.in({chany_top_in[61], chany_top_in[187], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size3 mux_right_track_96 (
		.in({chany_top_in[62], chany_top_in[191], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size3 mux_right_track_98 (
		.in({chany_top_in[64], chany_top_in[195], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size3 mux_right_track_100 (
		.in({chany_top_in[65], chany_top_in[199], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size3 mux_right_track_102 (
		.in({chany_top_in[66], chany_top_in[203], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size3 mux_right_track_104 (
		.in({chany_top_in[68], chany_top_in[207], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size3 mux_right_track_106 (
		.in({chany_top_in[69], chany_top_in[211], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size3 mux_right_track_108 (
		.in({chany_top_in[70], chany_top_in[215], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size3 mux_right_track_110 (
		.in({chany_top_in[72], chany_top_in[219], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size3 mux_right_track_112 (
		.in({chany_top_in[73], chany_top_in[223], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size3 mux_right_track_114 (
		.in({chany_top_in[74], chany_top_in[227], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size3 mux_right_track_116 (
		.in({chany_top_in[76], chany_top_in[231], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size3 mux_right_track_118 (
		.in({chany_top_in[77], chany_top_in[235], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size3 mux_right_track_120 (
		.in({chany_top_in[78], chany_top_in[239], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size3 mux_right_track_122 (
		.in({chany_top_in[80], chany_top_in[243], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_60_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size3 mux_right_track_124 (
		.in({chany_top_in[81], chany_top_in[247], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_61_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size3 mux_right_track_126 (
		.in({chany_top_in[82], chany_top_in[251], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_62_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size3 mux_right_track_128 (
		.in({chany_top_in[84], chany_top_in[255], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_63_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size3 mux_right_track_130 (
		.in({chany_top_in[85], chany_top_in[259], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_64_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size3 mux_right_track_132 (
		.in({chany_top_in[86], chany_top_in[263], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_65_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size3 mux_right_track_134 (
		.in({chany_top_in[88], chany_top_in[267], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_66_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size3 mux_right_track_136 (
		.in({chany_top_in[89], chany_top_in[271], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_67_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size3 mux_right_track_138 (
		.in({chany_top_in[90], chany_top_in[275], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_68_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size3 mux_right_track_140 (
		.in({chany_top_in[92], chany_top_in[279], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_69_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size3 mux_right_track_142 (
		.in({chany_top_in[93], chany_top_in[283], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_70_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size3 mux_right_track_144 (
		.in({chany_top_in[94], chany_top_in[287], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_71_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size3 mux_right_track_150 (
		.in({chany_top_in[98], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[292]}),
		.sram(mux_tree_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_72_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_size3 mux_right_track_152 (
		.in({chany_top_in[100], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[290]}),
		.sram(mux_tree_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_73_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size3 mux_right_track_154 (
		.in({chany_top_in[101], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[289]}),
		.sram(mux_tree_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_74_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_tree_tapbuf_size3 mux_right_track_156 (
		.in({chany_top_in[102], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[288]}),
		.sram(mux_tree_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_75_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_tree_tapbuf_size3 mux_right_track_158 (
		.in({chany_top_in[104], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[286]}),
		.sram(mux_tree_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_76_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_size3 mux_right_track_160 (
		.in({chany_top_in[105], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[285]}),
		.sram(mux_tree_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_77_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size3 mux_right_track_162 (
		.in({chany_top_in[106], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[284]}),
		.sram(mux_tree_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_78_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_tree_tapbuf_size3 mux_right_track_164 (
		.in({chany_top_in[108], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[282]}),
		.sram(mux_tree_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_79_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_tree_tapbuf_size3 mux_right_track_166 (
		.in({chany_top_in[109], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[281]}),
		.sram(mux_tree_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_80_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_size3 mux_right_track_168 (
		.in({chany_top_in[110], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[280]}),
		.sram(mux_tree_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_81_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size3 mux_right_track_170 (
		.in({chany_top_in[112], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[278]}),
		.sram(mux_tree_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_82_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_tree_tapbuf_size3 mux_right_track_172 (
		.in({chany_top_in[113], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[277]}),
		.sram(mux_tree_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_83_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_tree_tapbuf_size3 mux_right_track_174 (
		.in({chany_top_in[114], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[276]}),
		.sram(mux_tree_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_84_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_size3 mux_right_track_176 (
		.in({chany_top_in[116], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[274]}),
		.sram(mux_tree_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_85_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size3 mux_right_track_178 (
		.in({chany_top_in[117], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[273]}),
		.sram(mux_tree_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_tree_tapbuf_size3 mux_right_track_180 (
		.in({chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[272]}),
		.sram(mux_tree_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_tree_tapbuf_size3 mux_right_track_182 (
		.in({chany_top_in[120], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[270]}),
		.sram(mux_tree_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_size3 mux_right_track_184 (
		.in({chany_top_in[121], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[269]}),
		.sram(mux_tree_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_89_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size3 mux_right_track_186 (
		.in({chany_top_in[122], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[268]}),
		.sram(mux_tree_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_90_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_tree_tapbuf_size3 mux_right_track_188 (
		.in({chany_top_in[124], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[266]}),
		.sram(mux_tree_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_91_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_tree_tapbuf_size3 mux_right_track_190 (
		.in({chany_top_in[125], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[265]}),
		.sram(mux_tree_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_92_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_size3 mux_right_track_192 (
		.in({chany_top_in[126], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[264]}),
		.sram(mux_tree_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_93_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size3 mux_right_track_194 (
		.in({chany_top_in[128], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[262]}),
		.sram(mux_tree_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_94_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_tree_tapbuf_size3 mux_right_track_196 (
		.in({chany_top_in[129], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[261]}),
		.sram(mux_tree_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_95_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_tree_tapbuf_size3 mux_right_track_198 (
		.in({chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[260]}),
		.sram(mux_tree_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_96_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_tree_tapbuf_size3 mux_right_track_200 (
		.in({chany_top_in[132], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[258]}),
		.sram(mux_tree_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_97_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size3 mux_right_track_202 (
		.in({chany_top_in[133], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[257]}),
		.sram(mux_tree_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_98_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_tree_tapbuf_size3 mux_right_track_204 (
		.in({chany_top_in[134], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[256]}),
		.sram(mux_tree_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_99_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_tree_tapbuf_size3 mux_right_track_206 (
		.in({chany_top_in[136], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[254]}),
		.sram(mux_tree_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_100_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_tree_tapbuf_size3 mux_right_track_208 (
		.in({chany_top_in[137], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[253]}),
		.sram(mux_tree_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_101_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size3 mux_right_track_210 (
		.in({chany_top_in[138], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[252]}),
		.sram(mux_tree_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_102_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_tree_tapbuf_size3 mux_right_track_212 (
		.in({chany_top_in[140], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[250]}),
		.sram(mux_tree_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_103_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_tree_tapbuf_size3 mux_right_track_214 (
		.in({chany_top_in[141], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[249]}),
		.sram(mux_tree_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_104_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_tree_tapbuf_size3 mux_right_track_216 (
		.in({chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[248]}),
		.sram(mux_tree_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_105_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size3 mux_right_track_218 (
		.in({chany_top_in[144], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[246]}),
		.sram(mux_tree_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_106_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_tree_tapbuf_size3 mux_right_track_220 (
		.in({chany_top_in[145], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[245]}),
		.sram(mux_tree_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_107_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_tree_tapbuf_size3 mux_right_track_222 (
		.in({chany_top_in[146], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[244]}),
		.sram(mux_tree_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_108_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_tree_tapbuf_size3 mux_right_track_224 (
		.in({chany_top_in[148], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[242]}),
		.sram(mux_tree_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_109_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size3 mux_right_track_226 (
		.in({chany_top_in[149], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[241]}),
		.sram(mux_tree_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_110_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_tree_tapbuf_size3 mux_right_track_228 (
		.in({chany_top_in[150], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[240]}),
		.sram(mux_tree_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_111_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_tree_tapbuf_size3 mux_right_track_230 (
		.in({chany_top_in[152], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[238]}),
		.sram(mux_tree_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_112_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_tree_tapbuf_size3 mux_right_track_232 (
		.in({chany_top_in[153], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[237]}),
		.sram(mux_tree_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_113_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size3 mux_right_track_234 (
		.in({chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[236]}),
		.sram(mux_tree_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_114_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_tree_tapbuf_size3 mux_right_track_236 (
		.in({chany_top_in[156], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[234]}),
		.sram(mux_tree_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_115_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_tree_tapbuf_size3 mux_right_track_238 (
		.in({chany_top_in[157], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[233]}),
		.sram(mux_tree_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_116_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_tree_tapbuf_size3 mux_right_track_240 (
		.in({chany_top_in[158], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[232]}),
		.sram(mux_tree_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_117_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size3 mux_right_track_242 (
		.in({chany_top_in[160], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[230]}),
		.sram(mux_tree_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_118_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_tree_tapbuf_size3 mux_right_track_244 (
		.in({chany_top_in[161], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[229]}),
		.sram(mux_tree_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_119_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_tree_tapbuf_size3 mux_right_track_246 (
		.in({chany_top_in[162], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[228]}),
		.sram(mux_tree_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_tree_tapbuf_size3 mux_right_track_248 (
		.in({chany_top_in[164], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[226]}),
		.sram(mux_tree_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size3 mux_right_track_250 (
		.in({chany_top_in[165], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[225]}),
		.sram(mux_tree_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_tree_tapbuf_size3 mux_right_track_252 (
		.in({chany_top_in[166], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[224]}),
		.sram(mux_tree_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_tree_tapbuf_size3 mux_right_track_254 (
		.in({chany_top_in[168], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[222]}),
		.sram(mux_tree_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_tree_tapbuf_size3 mux_right_track_256 (
		.in({chany_top_in[169], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[221]}),
		.sram(mux_tree_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size3 mux_right_track_258 (
		.in({chany_top_in[170], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[220]}),
		.sram(mux_tree_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_tree_tapbuf_size3 mux_right_track_260 (
		.in({chany_top_in[172], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[218]}),
		.sram(mux_tree_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_tree_tapbuf_size3 mux_right_track_262 (
		.in({chany_top_in[173], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[217]}),
		.sram(mux_tree_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_tree_tapbuf_size3 mux_right_track_264 (
		.in({chany_top_in[174], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[216]}),
		.sram(mux_tree_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size3 mux_right_track_266 (
		.in({chany_top_in[176], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[214]}),
		.sram(mux_tree_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_tree_tapbuf_size3 mux_right_track_268 (
		.in({chany_top_in[177], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[213]}),
		.sram(mux_tree_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_tree_tapbuf_size3 mux_right_track_270 (
		.in({chany_top_in[178], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[212]}),
		.sram(mux_tree_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_tree_tapbuf_size3 mux_right_track_272 (
		.in({chany_top_in[180], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[210]}),
		.sram(mux_tree_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size3 mux_right_track_274 (
		.in({chany_top_in[181], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[209]}),
		.sram(mux_tree_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_tree_tapbuf_size3 mux_right_track_276 (
		.in({chany_top_in[182], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[208]}),
		.sram(mux_tree_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_tree_tapbuf_size3 mux_right_track_278 (
		.in({chany_top_in[184], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[206]}),
		.sram(mux_tree_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_tree_tapbuf_size3 mux_right_track_280 (
		.in({chany_top_in[185], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[205]}),
		.sram(mux_tree_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_137_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size3 mux_right_track_282 (
		.in({chany_top_in[186], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[204]}),
		.sram(mux_tree_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_138_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_tree_tapbuf_size3 mux_right_track_284 (
		.in({chany_top_in[188], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[202]}),
		.sram(mux_tree_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_139_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_tree_tapbuf_size3 mux_right_track_286 (
		.in({chany_top_in[189], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[201]}),
		.sram(mux_tree_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_140_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_tree_tapbuf_size3 mux_right_track_288 (
		.in({chany_top_in[190], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[200]}),
		.sram(mux_tree_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_141_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size3 mux_right_track_290 (
		.in({chany_top_in[192], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[198]}),
		.sram(mux_tree_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_142_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_tree_tapbuf_size3 mux_right_track_292 (
		.in({chany_top_in[193], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[197]}),
		.sram(mux_tree_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_143_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_tree_tapbuf_size3 mux_right_track_294 (
		.in({chany_top_in[194], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[196]}),
		.sram(mux_tree_tapbuf_size3_144_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_144_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_tree_tapbuf_size3 mux_right_track_296 (
		.in({chany_top_in[196], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[194]}),
		.sram(mux_tree_tapbuf_size3_145_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_145_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size3 mux_right_track_298 (
		.in({chany_top_in[197], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[193]}),
		.sram(mux_tree_tapbuf_size3_146_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_146_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_tree_tapbuf_size3 mux_right_track_300 (
		.in({chany_top_in[198], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[192]}),
		.sram(mux_tree_tapbuf_size3_147_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_147_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_tree_tapbuf_size3 mux_right_track_302 (
		.in({chany_top_in[200], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[190]}),
		.sram(mux_tree_tapbuf_size3_148_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_148_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_tree_tapbuf_size3 mux_right_track_304 (
		.in({chany_top_in[201], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[189]}),
		.sram(mux_tree_tapbuf_size3_149_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_149_sram_inv[0:1]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size3 mux_right_track_306 (
		.in({chany_top_in[202], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[188]}),
		.sram(mux_tree_tapbuf_size3_150_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_150_sram_inv[0:1]),
		.out(chanx_right_out[153]));

	mux_tree_tapbuf_size3 mux_right_track_308 (
		.in({chany_top_in[204], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[186]}),
		.sram(mux_tree_tapbuf_size3_151_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_151_sram_inv[0:1]),
		.out(chanx_right_out[154]));

	mux_tree_tapbuf_size3 mux_right_track_310 (
		.in({chany_top_in[205], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[185]}),
		.sram(mux_tree_tapbuf_size3_152_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_152_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_tree_tapbuf_size3 mux_right_track_312 (
		.in({chany_top_in[206], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[184]}),
		.sram(mux_tree_tapbuf_size3_153_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_153_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size3 mux_right_track_314 (
		.in({chany_top_in[208], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[182]}),
		.sram(mux_tree_tapbuf_size3_154_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_154_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_tree_tapbuf_size3 mux_right_track_316 (
		.in({chany_top_in[209], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[181]}),
		.sram(mux_tree_tapbuf_size3_155_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_155_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_tree_tapbuf_size3 mux_right_track_318 (
		.in({chany_top_in[210], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[180]}),
		.sram(mux_tree_tapbuf_size3_156_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_156_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_tree_tapbuf_size3 mux_right_track_320 (
		.in({chany_top_in[212], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[178]}),
		.sram(mux_tree_tapbuf_size3_157_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_157_sram_inv[0:1]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size3 mux_right_track_322 (
		.in({chany_top_in[213], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[177]}),
		.sram(mux_tree_tapbuf_size3_158_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_158_sram_inv[0:1]),
		.out(chanx_right_out[161]));

	mux_tree_tapbuf_size3 mux_right_track_324 (
		.in({chany_top_in[214], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[176]}),
		.sram(mux_tree_tapbuf_size3_159_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_159_sram_inv[0:1]),
		.out(chanx_right_out[162]));

	mux_tree_tapbuf_size3 mux_right_track_326 (
		.in({chany_top_in[216], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[174]}),
		.sram(mux_tree_tapbuf_size3_160_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_160_sram_inv[0:1]),
		.out(chanx_right_out[163]));

	mux_tree_tapbuf_size3 mux_right_track_328 (
		.in({chany_top_in[217], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[173]}),
		.sram(mux_tree_tapbuf_size3_161_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_161_sram_inv[0:1]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size3 mux_right_track_330 (
		.in({chany_top_in[218], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[172]}),
		.sram(mux_tree_tapbuf_size3_162_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_162_sram_inv[0:1]),
		.out(chanx_right_out[165]));

	mux_tree_tapbuf_size3 mux_right_track_332 (
		.in({chany_top_in[220], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[170]}),
		.sram(mux_tree_tapbuf_size3_163_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_163_sram_inv[0:1]),
		.out(chanx_right_out[166]));

	mux_tree_tapbuf_size3 mux_right_track_334 (
		.in({chany_top_in[221], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[169]}),
		.sram(mux_tree_tapbuf_size3_164_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_164_sram_inv[0:1]),
		.out(chanx_right_out[167]));

	mux_tree_tapbuf_size3 mux_right_track_336 (
		.in({chany_top_in[222], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[168]}),
		.sram(mux_tree_tapbuf_size3_165_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_165_sram_inv[0:1]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size3 mux_right_track_338 (
		.in({chany_top_in[224], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[166]}),
		.sram(mux_tree_tapbuf_size3_166_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_166_sram_inv[0:1]),
		.out(chanx_right_out[169]));

	mux_tree_tapbuf_size3 mux_right_track_340 (
		.in({chany_top_in[225], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[165]}),
		.sram(mux_tree_tapbuf_size3_167_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_167_sram_inv[0:1]),
		.out(chanx_right_out[170]));

	mux_tree_tapbuf_size3 mux_right_track_342 (
		.in({chany_top_in[226], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[164]}),
		.sram(mux_tree_tapbuf_size3_168_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_168_sram_inv[0:1]),
		.out(chanx_right_out[171]));

	mux_tree_tapbuf_size3 mux_right_track_344 (
		.in({chany_top_in[228], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[162]}),
		.sram(mux_tree_tapbuf_size3_169_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_169_sram_inv[0:1]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size3 mux_right_track_346 (
		.in({chany_top_in[229], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[161]}),
		.sram(mux_tree_tapbuf_size3_170_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_170_sram_inv[0:1]),
		.out(chanx_right_out[173]));

	mux_tree_tapbuf_size3 mux_right_track_348 (
		.in({chany_top_in[230], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[160]}),
		.sram(mux_tree_tapbuf_size3_171_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_171_sram_inv[0:1]),
		.out(chanx_right_out[174]));

	mux_tree_tapbuf_size3 mux_right_track_350 (
		.in({chany_top_in[232], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[158]}),
		.sram(mux_tree_tapbuf_size3_172_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_172_sram_inv[0:1]),
		.out(chanx_right_out[175]));

	mux_tree_tapbuf_size3 mux_right_track_352 (
		.in({chany_top_in[233], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[157]}),
		.sram(mux_tree_tapbuf_size3_173_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_173_sram_inv[0:1]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size3 mux_right_track_354 (
		.in({chany_top_in[234], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[156]}),
		.sram(mux_tree_tapbuf_size3_174_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_174_sram_inv[0:1]),
		.out(chanx_right_out[177]));

	mux_tree_tapbuf_size3 mux_right_track_356 (
		.in({chany_top_in[236], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[154]}),
		.sram(mux_tree_tapbuf_size3_175_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_175_sram_inv[0:1]),
		.out(chanx_right_out[178]));

	mux_tree_tapbuf_size3 mux_right_track_358 (
		.in({chany_top_in[237], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[153]}),
		.sram(mux_tree_tapbuf_size3_176_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_176_sram_inv[0:1]),
		.out(chanx_right_out[179]));

	mux_tree_tapbuf_size3 mux_right_track_360 (
		.in({chany_top_in[238], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[152]}),
		.sram(mux_tree_tapbuf_size3_177_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_177_sram_inv[0:1]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size3 mux_right_track_362 (
		.in({chany_top_in[240], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[150]}),
		.sram(mux_tree_tapbuf_size3_178_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_178_sram_inv[0:1]),
		.out(chanx_right_out[181]));

	mux_tree_tapbuf_size3 mux_right_track_364 (
		.in({chany_top_in[241], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[149]}),
		.sram(mux_tree_tapbuf_size3_179_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_179_sram_inv[0:1]),
		.out(chanx_right_out[182]));

	mux_tree_tapbuf_size3 mux_right_track_366 (
		.in({chany_top_in[242], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[148]}),
		.sram(mux_tree_tapbuf_size3_180_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_180_sram_inv[0:1]),
		.out(chanx_right_out[183]));

	mux_tree_tapbuf_size3 mux_right_track_368 (
		.in({chany_top_in[244], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[146]}),
		.sram(mux_tree_tapbuf_size3_181_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_181_sram_inv[0:1]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size3 mux_right_track_370 (
		.in({chany_top_in[245], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[145]}),
		.sram(mux_tree_tapbuf_size3_182_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_182_sram_inv[0:1]),
		.out(chanx_right_out[185]));

	mux_tree_tapbuf_size3 mux_right_track_372 (
		.in({chany_top_in[246], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[144]}),
		.sram(mux_tree_tapbuf_size3_183_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_183_sram_inv[0:1]),
		.out(chanx_right_out[186]));

	mux_tree_tapbuf_size3 mux_right_track_374 (
		.in({chany_top_in[248], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[142]}),
		.sram(mux_tree_tapbuf_size3_184_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_184_sram_inv[0:1]),
		.out(chanx_right_out[187]));

	mux_tree_tapbuf_size3 mux_right_track_376 (
		.in({chany_top_in[249], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[141]}),
		.sram(mux_tree_tapbuf_size3_185_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_185_sram_inv[0:1]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size3 mux_right_track_378 (
		.in({chany_top_in[250], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[140]}),
		.sram(mux_tree_tapbuf_size3_186_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_186_sram_inv[0:1]),
		.out(chanx_right_out[189]));

	mux_tree_tapbuf_size3 mux_right_track_380 (
		.in({chany_top_in[252], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[138]}),
		.sram(mux_tree_tapbuf_size3_187_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_187_sram_inv[0:1]),
		.out(chanx_right_out[190]));

	mux_tree_tapbuf_size3 mux_right_track_382 (
		.in({chany_top_in[253], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[137]}),
		.sram(mux_tree_tapbuf_size3_188_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_188_sram_inv[0:1]),
		.out(chanx_right_out[191]));

	mux_tree_tapbuf_size3 mux_right_track_384 (
		.in({chany_top_in[254], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[136]}),
		.sram(mux_tree_tapbuf_size3_189_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_189_sram_inv[0:1]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size3 mux_right_track_386 (
		.in({chany_top_in[256], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[134]}),
		.sram(mux_tree_tapbuf_size3_190_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_190_sram_inv[0:1]),
		.out(chanx_right_out[193]));

	mux_tree_tapbuf_size3 mux_right_track_388 (
		.in({chany_top_in[257], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[133]}),
		.sram(mux_tree_tapbuf_size3_191_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_191_sram_inv[0:1]),
		.out(chanx_right_out[194]));

	mux_tree_tapbuf_size3 mux_right_track_390 (
		.in({chany_top_in[258], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[132]}),
		.sram(mux_tree_tapbuf_size3_192_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_192_sram_inv[0:1]),
		.out(chanx_right_out[195]));

	mux_tree_tapbuf_size3 mux_right_track_392 (
		.in({chany_top_in[260], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[130]}),
		.sram(mux_tree_tapbuf_size3_193_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_193_sram_inv[0:1]),
		.out(chanx_right_out[196]));

	mux_tree_tapbuf_size3 mux_right_track_394 (
		.in({chany_top_in[261], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[129]}),
		.sram(mux_tree_tapbuf_size3_194_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_194_sram_inv[0:1]),
		.out(chanx_right_out[197]));

	mux_tree_tapbuf_size3 mux_right_track_396 (
		.in({chany_top_in[262], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[128]}),
		.sram(mux_tree_tapbuf_size3_195_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_195_sram_inv[0:1]),
		.out(chanx_right_out[198]));

	mux_tree_tapbuf_size3 mux_right_track_398 (
		.in({chany_top_in[264], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[126]}),
		.sram(mux_tree_tapbuf_size3_196_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_196_sram_inv[0:1]),
		.out(chanx_right_out[199]));

	mux_tree_tapbuf_size3 mux_right_track_400 (
		.in({chany_top_in[265], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[125]}),
		.sram(mux_tree_tapbuf_size3_197_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_197_sram_inv[0:1]),
		.out(chanx_right_out[200]));

	mux_tree_tapbuf_size3 mux_right_track_402 (
		.in({chany_top_in[266], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[124]}),
		.sram(mux_tree_tapbuf_size3_198_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_198_sram_inv[0:1]),
		.out(chanx_right_out[201]));

	mux_tree_tapbuf_size3 mux_right_track_404 (
		.in({chany_top_in[268], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[122]}),
		.sram(mux_tree_tapbuf_size3_199_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_199_sram_inv[0:1]),
		.out(chanx_right_out[202]));

	mux_tree_tapbuf_size3 mux_right_track_406 (
		.in({chany_top_in[269], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[121]}),
		.sram(mux_tree_tapbuf_size3_200_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_200_sram_inv[0:1]),
		.out(chanx_right_out[203]));

	mux_tree_tapbuf_size3 mux_right_track_408 (
		.in({chany_top_in[270], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[120]}),
		.sram(mux_tree_tapbuf_size3_201_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_201_sram_inv[0:1]),
		.out(chanx_right_out[204]));

	mux_tree_tapbuf_size3 mux_right_track_410 (
		.in({chany_top_in[272], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[118]}),
		.sram(mux_tree_tapbuf_size3_202_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_202_sram_inv[0:1]),
		.out(chanx_right_out[205]));

	mux_tree_tapbuf_size3 mux_right_track_412 (
		.in({chany_top_in[273], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[117]}),
		.sram(mux_tree_tapbuf_size3_203_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_203_sram_inv[0:1]),
		.out(chanx_right_out[206]));

	mux_tree_tapbuf_size3 mux_right_track_414 (
		.in({chany_top_in[274], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[116]}),
		.sram(mux_tree_tapbuf_size3_204_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_204_sram_inv[0:1]),
		.out(chanx_right_out[207]));

	mux_tree_tapbuf_size3 mux_right_track_416 (
		.in({chany_top_in[276], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[114]}),
		.sram(mux_tree_tapbuf_size3_205_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_205_sram_inv[0:1]),
		.out(chanx_right_out[208]));

	mux_tree_tapbuf_size3 mux_right_track_418 (
		.in({chany_top_in[277], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[113]}),
		.sram(mux_tree_tapbuf_size3_206_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_206_sram_inv[0:1]),
		.out(chanx_right_out[209]));

	mux_tree_tapbuf_size3 mux_right_track_420 (
		.in({chany_top_in[278], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[112]}),
		.sram(mux_tree_tapbuf_size3_207_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_207_sram_inv[0:1]),
		.out(chanx_right_out[210]));

	mux_tree_tapbuf_size3 mux_right_track_422 (
		.in({chany_top_in[280], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[110]}),
		.sram(mux_tree_tapbuf_size3_208_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_208_sram_inv[0:1]),
		.out(chanx_right_out[211]));

	mux_tree_tapbuf_size3 mux_right_track_424 (
		.in({chany_top_in[281], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[109]}),
		.sram(mux_tree_tapbuf_size3_209_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_209_sram_inv[0:1]),
		.out(chanx_right_out[212]));

	mux_tree_tapbuf_size3 mux_right_track_426 (
		.in({chany_top_in[282], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[108]}),
		.sram(mux_tree_tapbuf_size3_210_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_210_sram_inv[0:1]),
		.out(chanx_right_out[213]));

	mux_tree_tapbuf_size3 mux_right_track_428 (
		.in({chany_top_in[284], right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[106]}),
		.sram(mux_tree_tapbuf_size3_211_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_211_sram_inv[0:1]),
		.out(chanx_right_out[214]));

	mux_tree_tapbuf_size3 mux_right_track_430 (
		.in({chany_top_in[285], right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[105]}),
		.sram(mux_tree_tapbuf_size3_212_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_212_sram_inv[0:1]),
		.out(chanx_right_out[215]));

	mux_tree_tapbuf_size3 mux_right_track_432 (
		.in({chany_top_in[286], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[104]}),
		.sram(mux_tree_tapbuf_size3_213_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_213_sram_inv[0:1]),
		.out(chanx_right_out[216]));

	mux_tree_tapbuf_size3 mux_right_track_434 (
		.in({chany_top_in[288], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size3_214_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_214_sram_inv[0:1]),
		.out(chanx_right_out[217]));

	mux_tree_tapbuf_size3 mux_right_track_436 (
		.in({chany_top_in[289], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size3_215_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_215_sram_inv[0:1]),
		.out(chanx_right_out[218]));

	mux_tree_tapbuf_size3 mux_right_track_438 (
		.in({chany_top_in[290], right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size3_216_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_216_sram_inv[0:1]),
		.out(chanx_right_out[219]));

	mux_tree_tapbuf_size3 mux_right_track_440 (
		.in({chany_top_in[292], right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size3_217_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_217_sram_inv[0:1]),
		.out(chanx_right_out[220]));

	mux_tree_tapbuf_size3 mux_right_track_446 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[94], chany_bottom_in[287]}),
		.sram(mux_tree_tapbuf_size3_218_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_218_sram_inv[0:1]),
		.out(chanx_right_out[223]));

	mux_tree_tapbuf_size3 mux_right_track_448 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[93], chany_bottom_in[283]}),
		.sram(mux_tree_tapbuf_size3_219_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_219_sram_inv[0:1]),
		.out(chanx_right_out[224]));

	mux_tree_tapbuf_size3 mux_right_track_450 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[92], chany_bottom_in[279]}),
		.sram(mux_tree_tapbuf_size3_220_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_220_sram_inv[0:1]),
		.out(chanx_right_out[225]));

	mux_tree_tapbuf_size3 mux_right_track_452 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[90], chany_bottom_in[275]}),
		.sram(mux_tree_tapbuf_size3_221_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_221_sram_inv[0:1]),
		.out(chanx_right_out[226]));

	mux_tree_tapbuf_size3 mux_right_track_454 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[89], chany_bottom_in[271]}),
		.sram(mux_tree_tapbuf_size3_222_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_222_sram_inv[0:1]),
		.out(chanx_right_out[227]));

	mux_tree_tapbuf_size3 mux_right_track_456 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[88], chany_bottom_in[267]}),
		.sram(mux_tree_tapbuf_size3_223_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_223_sram_inv[0:1]),
		.out(chanx_right_out[228]));

	mux_tree_tapbuf_size3 mux_right_track_458 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[86], chany_bottom_in[263]}),
		.sram(mux_tree_tapbuf_size3_224_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_224_sram_inv[0:1]),
		.out(chanx_right_out[229]));

	mux_tree_tapbuf_size3 mux_right_track_460 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[85], chany_bottom_in[259]}),
		.sram(mux_tree_tapbuf_size3_225_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_225_sram_inv[0:1]),
		.out(chanx_right_out[230]));

	mux_tree_tapbuf_size3 mux_right_track_462 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[84], chany_bottom_in[255]}),
		.sram(mux_tree_tapbuf_size3_226_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_226_sram_inv[0:1]),
		.out(chanx_right_out[231]));

	mux_tree_tapbuf_size3 mux_right_track_464 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[82], chany_bottom_in[251]}),
		.sram(mux_tree_tapbuf_size3_227_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_227_sram_inv[0:1]),
		.out(chanx_right_out[232]));

	mux_tree_tapbuf_size3 mux_right_track_466 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[81], chany_bottom_in[247]}),
		.sram(mux_tree_tapbuf_size3_228_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_228_sram_inv[0:1]),
		.out(chanx_right_out[233]));

	mux_tree_tapbuf_size3 mux_right_track_468 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[80], chany_bottom_in[243]}),
		.sram(mux_tree_tapbuf_size3_229_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_229_sram_inv[0:1]),
		.out(chanx_right_out[234]));

	mux_tree_tapbuf_size3 mux_right_track_470 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[78], chany_bottom_in[239]}),
		.sram(mux_tree_tapbuf_size3_230_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_230_sram_inv[0:1]),
		.out(chanx_right_out[235]));

	mux_tree_tapbuf_size3 mux_right_track_472 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[77], chany_bottom_in[235]}),
		.sram(mux_tree_tapbuf_size3_231_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_231_sram_inv[0:1]),
		.out(chanx_right_out[236]));

	mux_tree_tapbuf_size3 mux_right_track_474 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[76], chany_bottom_in[231]}),
		.sram(mux_tree_tapbuf_size3_232_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_232_sram_inv[0:1]),
		.out(chanx_right_out[237]));

	mux_tree_tapbuf_size3 mux_right_track_476 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[74], chany_bottom_in[227]}),
		.sram(mux_tree_tapbuf_size3_233_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_233_sram_inv[0:1]),
		.out(chanx_right_out[238]));

	mux_tree_tapbuf_size3 mux_right_track_478 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[73], chany_bottom_in[223]}),
		.sram(mux_tree_tapbuf_size3_234_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_234_sram_inv[0:1]),
		.out(chanx_right_out[239]));

	mux_tree_tapbuf_size3 mux_right_track_480 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[72], chany_bottom_in[219]}),
		.sram(mux_tree_tapbuf_size3_235_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_235_sram_inv[0:1]),
		.out(chanx_right_out[240]));

	mux_tree_tapbuf_size3 mux_right_track_482 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[70], chany_bottom_in[215]}),
		.sram(mux_tree_tapbuf_size3_236_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_236_sram_inv[0:1]),
		.out(chanx_right_out[241]));

	mux_tree_tapbuf_size3 mux_right_track_484 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[69], chany_bottom_in[211]}),
		.sram(mux_tree_tapbuf_size3_237_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_237_sram_inv[0:1]),
		.out(chanx_right_out[242]));

	mux_tree_tapbuf_size3 mux_right_track_486 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[68], chany_bottom_in[207]}),
		.sram(mux_tree_tapbuf_size3_238_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_238_sram_inv[0:1]),
		.out(chanx_right_out[243]));

	mux_tree_tapbuf_size3 mux_right_track_488 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[66], chany_bottom_in[203]}),
		.sram(mux_tree_tapbuf_size3_239_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_239_sram_inv[0:1]),
		.out(chanx_right_out[244]));

	mux_tree_tapbuf_size3 mux_right_track_490 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[65], chany_bottom_in[199]}),
		.sram(mux_tree_tapbuf_size3_240_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_240_sram_inv[0:1]),
		.out(chanx_right_out[245]));

	mux_tree_tapbuf_size3 mux_right_track_492 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[64], chany_bottom_in[195]}),
		.sram(mux_tree_tapbuf_size3_241_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_241_sram_inv[0:1]),
		.out(chanx_right_out[246]));

	mux_tree_tapbuf_size3 mux_right_track_494 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[62], chany_bottom_in[191]}),
		.sram(mux_tree_tapbuf_size3_242_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_242_sram_inv[0:1]),
		.out(chanx_right_out[247]));

	mux_tree_tapbuf_size3 mux_right_track_496 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[61], chany_bottom_in[187]}),
		.sram(mux_tree_tapbuf_size3_243_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_243_sram_inv[0:1]),
		.out(chanx_right_out[248]));

	mux_tree_tapbuf_size3 mux_right_track_498 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[60], chany_bottom_in[183]}),
		.sram(mux_tree_tapbuf_size3_244_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_244_sram_inv[0:1]),
		.out(chanx_right_out[249]));

	mux_tree_tapbuf_size3 mux_right_track_500 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[58], chany_bottom_in[179]}),
		.sram(mux_tree_tapbuf_size3_245_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_245_sram_inv[0:1]),
		.out(chanx_right_out[250]));

	mux_tree_tapbuf_size3 mux_right_track_502 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[57], chany_bottom_in[175]}),
		.sram(mux_tree_tapbuf_size3_246_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_246_sram_inv[0:1]),
		.out(chanx_right_out[251]));

	mux_tree_tapbuf_size3 mux_right_track_504 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[56], chany_bottom_in[171]}),
		.sram(mux_tree_tapbuf_size3_247_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_247_sram_inv[0:1]),
		.out(chanx_right_out[252]));

	mux_tree_tapbuf_size3 mux_right_track_506 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[54], chany_bottom_in[167]}),
		.sram(mux_tree_tapbuf_size3_248_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_248_sram_inv[0:1]),
		.out(chanx_right_out[253]));

	mux_tree_tapbuf_size3 mux_right_track_508 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[53], chany_bottom_in[163]}),
		.sram(mux_tree_tapbuf_size3_249_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_249_sram_inv[0:1]),
		.out(chanx_right_out[254]));

	mux_tree_tapbuf_size3 mux_right_track_510 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[52], chany_bottom_in[159]}),
		.sram(mux_tree_tapbuf_size3_250_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_250_sram_inv[0:1]),
		.out(chanx_right_out[255]));

	mux_tree_tapbuf_size3 mux_right_track_512 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[50], chany_bottom_in[155]}),
		.sram(mux_tree_tapbuf_size3_251_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_251_sram_inv[0:1]),
		.out(chanx_right_out[256]));

	mux_tree_tapbuf_size3 mux_right_track_514 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[49], chany_bottom_in[151]}),
		.sram(mux_tree_tapbuf_size3_252_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_252_sram_inv[0:1]),
		.out(chanx_right_out[257]));

	mux_tree_tapbuf_size3 mux_right_track_516 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[48], chany_bottom_in[147]}),
		.sram(mux_tree_tapbuf_size3_253_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_253_sram_inv[0:1]),
		.out(chanx_right_out[258]));

	mux_tree_tapbuf_size3 mux_right_track_518 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[46], chany_bottom_in[143]}),
		.sram(mux_tree_tapbuf_size3_254_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_254_sram_inv[0:1]),
		.out(chanx_right_out[259]));

	mux_tree_tapbuf_size3 mux_right_track_520 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[45], chany_bottom_in[139]}),
		.sram(mux_tree_tapbuf_size3_255_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_255_sram_inv[0:1]),
		.out(chanx_right_out[260]));

	mux_tree_tapbuf_size3 mux_right_track_522 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[44], chany_bottom_in[135]}),
		.sram(mux_tree_tapbuf_size3_256_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_256_sram_inv[0:1]),
		.out(chanx_right_out[261]));

	mux_tree_tapbuf_size3 mux_right_track_524 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[42], chany_bottom_in[131]}),
		.sram(mux_tree_tapbuf_size3_257_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_257_sram_inv[0:1]),
		.out(chanx_right_out[262]));

	mux_tree_tapbuf_size3 mux_right_track_526 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[41], chany_bottom_in[127]}),
		.sram(mux_tree_tapbuf_size3_258_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_258_sram_inv[0:1]),
		.out(chanx_right_out[263]));

	mux_tree_tapbuf_size3 mux_right_track_528 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[40], chany_bottom_in[123]}),
		.sram(mux_tree_tapbuf_size3_259_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_259_sram_inv[0:1]),
		.out(chanx_right_out[264]));

	mux_tree_tapbuf_size3 mux_right_track_530 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[38], chany_bottom_in[119]}),
		.sram(mux_tree_tapbuf_size3_260_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_260_sram_inv[0:1]),
		.out(chanx_right_out[265]));

	mux_tree_tapbuf_size3 mux_right_track_532 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[37], chany_bottom_in[115]}),
		.sram(mux_tree_tapbuf_size3_261_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_261_sram_inv[0:1]),
		.out(chanx_right_out[266]));

	mux_tree_tapbuf_size3 mux_right_track_534 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[36], chany_bottom_in[111]}),
		.sram(mux_tree_tapbuf_size3_262_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_262_sram_inv[0:1]),
		.out(chanx_right_out[267]));

	mux_tree_tapbuf_size3 mux_right_track_536 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[34], chany_bottom_in[107]}),
		.sram(mux_tree_tapbuf_size3_263_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_263_sram_inv[0:1]),
		.out(chanx_right_out[268]));

	mux_tree_tapbuf_size3 mux_right_track_538 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[33], chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size3_264_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_264_sram_inv[0:1]),
		.out(chanx_right_out[269]));

	mux_tree_tapbuf_size3 mux_right_track_540 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[32], chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size3_265_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_265_sram_inv[0:1]),
		.out(chanx_right_out[270]));

	mux_tree_tapbuf_size3 mux_right_track_542 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[30], chany_bottom_in[95]}),
		.sram(mux_tree_tapbuf_size3_266_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_266_sram_inv[0:1]),
		.out(chanx_right_out[271]));

	mux_tree_tapbuf_size3 mux_right_track_544 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[29], chany_bottom_in[91]}),
		.sram(mux_tree_tapbuf_size3_267_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_267_sram_inv[0:1]),
		.out(chanx_right_out[272]));

	mux_tree_tapbuf_size3 mux_right_track_546 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[28], chany_bottom_in[87]}),
		.sram(mux_tree_tapbuf_size3_268_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_268_sram_inv[0:1]),
		.out(chanx_right_out[273]));

	mux_tree_tapbuf_size3 mux_right_track_548 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[26], chany_bottom_in[83]}),
		.sram(mux_tree_tapbuf_size3_269_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_269_sram_inv[0:1]),
		.out(chanx_right_out[274]));

	mux_tree_tapbuf_size3 mux_right_track_550 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[25], chany_bottom_in[79]}),
		.sram(mux_tree_tapbuf_size3_270_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_270_sram_inv[0:1]),
		.out(chanx_right_out[275]));

	mux_tree_tapbuf_size3 mux_right_track_552 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_size3_271_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_271_sram_inv[0:1]),
		.out(chanx_right_out[276]));

	mux_tree_tapbuf_size3 mux_right_track_554 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_size3_272_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_272_sram_inv[0:1]),
		.out(chanx_right_out[277]));

	mux_tree_tapbuf_size3 mux_right_track_556 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size3_273_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_273_sram_inv[0:1]),
		.out(chanx_right_out[278]));

	mux_tree_tapbuf_size3 mux_right_track_558 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size3_274_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_274_sram_inv[0:1]),
		.out(chanx_right_out[279]));

	mux_tree_tapbuf_size3 mux_right_track_560 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size3_275_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_275_sram_inv[0:1]),
		.out(chanx_right_out[280]));

	mux_tree_tapbuf_size3 mux_right_track_562 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size3_276_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_276_sram_inv[0:1]),
		.out(chanx_right_out[281]));

	mux_tree_tapbuf_size3 mux_right_track_564 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size3_277_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_277_sram_inv[0:1]),
		.out(chanx_right_out[282]));

	mux_tree_tapbuf_size3 mux_right_track_566 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size3_278_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_278_sram_inv[0:1]),
		.out(chanx_right_out[283]));

	mux_tree_tapbuf_size3 mux_right_track_568 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size3_279_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_279_sram_inv[0:1]),
		.out(chanx_right_out[284]));

	mux_tree_tapbuf_size3 mux_right_track_570 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size3_280_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_280_sram_inv[0:1]),
		.out(chanx_right_out[285]));

	mux_tree_tapbuf_size3 mux_right_track_572 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size3_281_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_281_sram_inv[0:1]),
		.out(chanx_right_out[286]));

	mux_tree_tapbuf_size3 mux_right_track_574 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size3_282_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_282_sram_inv[0:1]),
		.out(chanx_right_out[287]));

	mux_tree_tapbuf_size3 mux_right_track_576 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size3_283_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_283_sram_inv[0:1]),
		.out(chanx_right_out[288]));

	mux_tree_tapbuf_size3 mux_right_track_578 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size3_284_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_284_sram_inv[0:1]),
		.out(chanx_right_out[289]));

	mux_tree_tapbuf_size3 mux_right_track_580 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size3_285_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_285_sram_inv[0:1]),
		.out(chanx_right_out[290]));

	mux_tree_tapbuf_size3 mux_right_track_582 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_, chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size3_286_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_286_sram_inv[0:1]),
		.out(chanx_right_out[291]));

	mux_tree_tapbuf_size3 mux_right_track_584 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size3_287_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_287_sram_inv[0:1]),
		.out(chanx_right_out[292]));

	mux_tree_tapbuf_size3 mux_right_track_586 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size3_288_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_288_sram_inv[0:1]),
		.out(chanx_right_out[293]));

	mux_tree_tapbuf_size3 mux_right_track_588 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_size3_289_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_289_sram_inv[0:1]),
		.out(chanx_right_out[294]));

	mux_tree_tapbuf_size3_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_60_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_61_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_62_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_63_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_64_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_65_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_66_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_67_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_68_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_69_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_70_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_71_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_72_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_73_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_74_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_75_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_76_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_77_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_78_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_79_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_80_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_81_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_82_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_83_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_84_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_85_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_86_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_87_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_88_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_89_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_90_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_91_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_92_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_93_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_94_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_95_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_96_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_97_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_98_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_99_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_100_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_101_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_102_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_103_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_104_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_105_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_106_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_107_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_108_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_109_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_110_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_111_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_112_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_113_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_114_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_115_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_116_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_117_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_118_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_119_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_120_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_121_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_122_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_123_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_124_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_125_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_126_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_127_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_128_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_129_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_130_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_131_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_132_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_133_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_134_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_135_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_136_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_137_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_138_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_139_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_140_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_141_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_142_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_143_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_144_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_144_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_145_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_145_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_146_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_146_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_147_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_147_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_148_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_148_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_149_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_149_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_150_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_150_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_151_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_151_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_152_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_152_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_153_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_153_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_154_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_154_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_155_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_155_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_156_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_156_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_157_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_157_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_158_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_158_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_159_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_159_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_160_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_160_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_161_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_161_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_162_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_162_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_163_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_163_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_164_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_164_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_165_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_165_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_166_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_166_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_167_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_167_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_168_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_168_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_169_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_169_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_170_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_170_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_171_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_171_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_172_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_172_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_173_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_173_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_174_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_174_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_175_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_175_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_176_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_176_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_177_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_177_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_178_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_178_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_179_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_179_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_180_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_180_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_181_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_181_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_182_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_182_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_183_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_183_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_184_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_184_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_185_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_185_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_378 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_186_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_186_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_380 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_187_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_187_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_382 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_188_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_188_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_189_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_189_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_386 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_190_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_190_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_388 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_191_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_191_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_390 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_192_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_192_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_193_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_193_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_394 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_194_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_194_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_396 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_195_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_195_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_398 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_196_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_196_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_197_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_197_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_402 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_198_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_198_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_404 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_199_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_199_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_406 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_200_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_200_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_201_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_201_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_410 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_202_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_202_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_412 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_203_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_203_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_414 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_204_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_204_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_205_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_205_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_418 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_206_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_206_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_420 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_207_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_207_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_422 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_208_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_208_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_209_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_209_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_426 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_210_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_210_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_428 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_211_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_211_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_430 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_212_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_212_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_213_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_213_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_434 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_214_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_214_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_436 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_215_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_215_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_438 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_216_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_216_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_217_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_217_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_446 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_218_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_218_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_219_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_219_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_450 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_220_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_220_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_452 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_221_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_221_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_454 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_222_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_222_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_223_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_223_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_458 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_224_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_224_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_460 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_224_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_225_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_225_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_225_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_462 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_225_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_226_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_226_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_226_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_226_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_227_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_227_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_227_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_466 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_227_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_228_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_228_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_228_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_468 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_228_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_229_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_229_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_229_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_470 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_229_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_230_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_230_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_230_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_230_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_231_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_231_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_231_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_474 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_231_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_232_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_232_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_232_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_476 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_232_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_233_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_233_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_233_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_478 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_233_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_234_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_234_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_234_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_234_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_235_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_235_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_235_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_482 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_235_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_236_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_236_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_236_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_484 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_236_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_237_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_237_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_237_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_486 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_237_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_238_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_238_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_238_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_238_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_239_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_239_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_239_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_490 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_239_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_240_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_240_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_240_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_492 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_240_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_241_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_241_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_241_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_494 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_241_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_242_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_242_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_242_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_242_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_243_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_243_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_243_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_498 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_243_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_244_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_244_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_244_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_500 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_244_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_245_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_245_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_245_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_502 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_245_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_246_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_246_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_246_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_246_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_247_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_247_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_247_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_506 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_247_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_248_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_248_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_248_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_508 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_248_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_249_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_249_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_249_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_510 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_249_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_250_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_250_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_250_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_250_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_251_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_251_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_251_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_514 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_251_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_252_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_252_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_252_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_516 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_252_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_253_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_253_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_253_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_518 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_253_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_254_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_254_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_254_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_254_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_255_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_255_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_255_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_522 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_255_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_256_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_256_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_256_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_524 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_256_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_257_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_257_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_257_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_526 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_257_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_258_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_258_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_258_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_258_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_259_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_259_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_259_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_530 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_259_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_260_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_260_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_260_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_532 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_260_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_261_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_261_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_261_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_534 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_261_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_262_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_262_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_262_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_262_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_263_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_263_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_263_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_538 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_263_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_264_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_264_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_264_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_540 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_264_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_265_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_265_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_265_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_542 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_265_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_266_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_266_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_266_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_266_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_267_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_267_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_267_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_546 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_267_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_268_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_268_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_268_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_548 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_268_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_269_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_269_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_269_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_550 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_269_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_270_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_270_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_270_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_270_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_271_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_271_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_271_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_554 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_271_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_272_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_272_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_272_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_556 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_272_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_273_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_273_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_273_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_558 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_273_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_274_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_274_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_274_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_274_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_275_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_275_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_275_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_562 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_275_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_276_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_276_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_276_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_564 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_276_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_277_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_277_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_277_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_566 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_277_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_278_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_278_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_278_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_278_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_279_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_279_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_279_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_570 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_279_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_280_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_280_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_280_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_572 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_280_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_281_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_281_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_281_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_574 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_281_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_282_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_282_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_282_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_576 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_282_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_283_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_283_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_283_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_578 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_283_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_284_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_284_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_284_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_580 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_284_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_285_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_285_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_285_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_582 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_285_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_286_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_286_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_286_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_584 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_286_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_287_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_287_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_287_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_586 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_287_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_288_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_288_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_288_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_588 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_288_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_289_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_289_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_289_sram_inv[0:1]));

	mux_tree_tapbuf_size4 mux_right_track_146 (
		.in({chany_top_in[96], chany_top_in[291], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, chany_bottom_in[294]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chanx_right_out[73]));

	mux_tree_tapbuf_size4 mux_right_track_148 (
		.in({chany_top_in[97], chany_top_in[295], right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, chany_bottom_in[293]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chanx_right_out[74]));

	mux_tree_tapbuf_size4 mux_right_track_442 (
		.in({chany_top_in[293], right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_, chany_bottom_in[97], chany_bottom_in[295]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chanx_right_out[221]));

	mux_tree_tapbuf_size4 mux_right_track_444 (
		.in({chany_top_in[294], right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_, chany_bottom_in[96], chany_bottom_in[291]}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chanx_right_out[222]));

	mux_tree_tapbuf_size4_mem mem_right_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_442 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_444 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7 mux_bottom_track_1 (
		.in({chanx_right_in[72], chanx_right_in[146], chanx_right_in[220], chanx_right_in[294], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size7 mux_bottom_track_9 (
		.in({chanx_right_in[71], chanx_right_in[145], chanx_right_in[219], chanx_right_in[293], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size7 mux_bottom_track_17 (
		.in({chanx_right_in[70], chanx_right_in[144], chanx_right_in[218], chanx_right_in[292], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size7 mux_bottom_track_25 (
		.in({chanx_right_in[69], chanx_right_in[143], chanx_right_in[217], chanx_right_in[291], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size7 mux_bottom_track_33 (
		.in({chanx_right_in[68], chanx_right_in[142], chanx_right_in[216], chanx_right_in[290], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_4_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size7 mux_bottom_track_73 (
		.in({chanx_right_in[63], chanx_right_in[137], chanx_right_in[211], chanx_right_in[285], bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_5_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size7 mux_bottom_track_81 (
		.in({chanx_right_in[62], chanx_right_in[136], chanx_right_in[210], chanx_right_in[284], bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_6_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size7 mux_bottom_track_89 (
		.in({chanx_right_in[61], chanx_right_in[135], chanx_right_in[209], chanx_right_in[283], bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_7_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size7 mux_bottom_track_97 (
		.in({chanx_right_in[60], chanx_right_in[134], chanx_right_in[208], chanx_right_in[282], bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_8_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size7 mux_bottom_track_105 (
		.in({chanx_right_in[59], chanx_right_in[133], chanx_right_in[207], chanx_right_in[281], bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_9_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_289_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_9_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_0__4_ -----

//----- Default net type -----
`default_nettype wire



