//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 12:51:27 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for fpga_top -----
module fpga_top(prog_clk,
                set,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:159] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__0_ccff_tail;
wire [0:192] cbx_1__0__0_chanx_left_out;
wire [0:192] cbx_1__0__0_chanx_right_out;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__1_ccff_tail;
wire [0:192] cbx_1__0__1_chanx_left_out;
wire [0:192] cbx_1__0__1_chanx_right_out;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__2_ccff_tail;
wire [0:192] cbx_1__0__2_chanx_left_out;
wire [0:192] cbx_1__0__2_chanx_right_out;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__0__3_ccff_tail;
wire [0:192] cbx_1__0__3_chanx_left_out;
wire [0:192] cbx_1__0__3_chanx_right_out;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__1__0_ccff_tail;
wire [0:192] cbx_1__1__0_chanx_left_out;
wire [0:192] cbx_1__1__0_chanx_right_out;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_;
wire [0:0] cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__1__1_ccff_tail;
wire [0:192] cbx_1__1__1_chanx_left_out;
wire [0:192] cbx_1__1__1_chanx_right_out;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_;
wire [0:0] cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__1__2_ccff_tail;
wire [0:192] cbx_1__1__2_chanx_left_out;
wire [0:192] cbx_1__1__2_chanx_right_out;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_;
wire [0:0] cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__1__3_ccff_tail;
wire [0:192] cbx_1__1__3_chanx_left_out;
wire [0:192] cbx_1__1__3_chanx_right_out;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_;
wire [0:0] cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_;
wire [0:0] cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_;
wire [0:0] cbx_1__2__0_ccff_tail;
wire [0:192] cbx_1__2__0_chanx_left_out;
wire [0:192] cbx_1__2__0_chanx_right_out;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_;
wire [0:0] cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_;
wire [0:0] cbx_1__2__1_ccff_tail;
wire [0:192] cbx_1__2__1_chanx_left_out;
wire [0:192] cbx_1__2__1_chanx_right_out;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_;
wire [0:0] cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_;
wire [0:0] cbx_1__2__2_ccff_tail;
wire [0:192] cbx_1__2__2_chanx_left_out;
wire [0:192] cbx_1__2__2_chanx_right_out;
wire [0:0] cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_;
wire [0:0] cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_;
wire [0:0] cbx_1__2__3_ccff_tail;
wire [0:192] cbx_1__2__3_chanx_left_out;
wire [0:192] cbx_1__2__3_chanx_right_out;
wire [0:0] cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__0_ccff_tail;
wire [0:192] cbx_1__3__0_chanx_left_out;
wire [0:192] cbx_1__3__0_chanx_right_out;
wire [0:0] cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__10_ccff_tail;
wire [0:192] cbx_1__3__10_chanx_left_out;
wire [0:192] cbx_1__3__10_chanx_right_out;
wire [0:0] cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__11_ccff_tail;
wire [0:192] cbx_1__3__11_chanx_left_out;
wire [0:192] cbx_1__3__11_chanx_right_out;
wire [0:0] cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__1_ccff_tail;
wire [0:192] cbx_1__3__1_chanx_left_out;
wire [0:192] cbx_1__3__1_chanx_right_out;
wire [0:0] cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__2_ccff_tail;
wire [0:192] cbx_1__3__2_chanx_left_out;
wire [0:192] cbx_1__3__2_chanx_right_out;
wire [0:0] cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__3_ccff_tail;
wire [0:192] cbx_1__3__3_chanx_left_out;
wire [0:192] cbx_1__3__3_chanx_right_out;
wire [0:0] cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__4_ccff_tail;
wire [0:192] cbx_1__3__4_chanx_left_out;
wire [0:192] cbx_1__3__4_chanx_right_out;
wire [0:0] cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__5_ccff_tail;
wire [0:192] cbx_1__3__5_chanx_left_out;
wire [0:192] cbx_1__3__5_chanx_right_out;
wire [0:0] cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__6_ccff_tail;
wire [0:192] cbx_1__3__6_chanx_left_out;
wire [0:192] cbx_1__3__6_chanx_right_out;
wire [0:0] cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__7_ccff_tail;
wire [0:192] cbx_1__3__7_chanx_left_out;
wire [0:192] cbx_1__3__7_chanx_right_out;
wire [0:0] cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__8_ccff_tail;
wire [0:192] cbx_1__3__8_chanx_left_out;
wire [0:192] cbx_1__3__8_chanx_right_out;
wire [0:0] cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__3__9_ccff_tail;
wire [0:192] cbx_1__3__9_chanx_left_out;
wire [0:192] cbx_1__3__9_chanx_right_out;
wire [0:0] cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_;
wire [0:0] cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_;
wire [0:0] cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__6__0_ccff_tail;
wire [0:192] cbx_1__6__0_chanx_left_out;
wire [0:192] cbx_1__6__0_chanx_right_out;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__6__1_ccff_tail;
wire [0:192] cbx_1__6__1_chanx_left_out;
wire [0:192] cbx_1__6__1_chanx_right_out;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__6__2_ccff_tail;
wire [0:192] cbx_1__6__2_chanx_left_out;
wire [0:192] cbx_1__6__2_chanx_right_out;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_;
wire [0:0] cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_;
wire [0:0] cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_;
wire [0:0] cbx_1__6__3_ccff_tail;
wire [0:192] cbx_1__6__3_chanx_left_out;
wire [0:192] cbx_1__6__3_chanx_right_out;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__0_ccff_tail;
wire [0:192] cby_0__1__0_chany_bottom_out;
wire [0:192] cby_0__1__0_chany_top_out;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__1__1_ccff_tail;
wire [0:192] cby_0__1__1_chany_bottom_out;
wire [0:192] cby_0__1__1_chany_top_out;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__1__2_ccff_tail;
wire [0:192] cby_0__1__2_chany_bottom_out;
wire [0:192] cby_0__1__2_chany_top_out;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__1__3_ccff_tail;
wire [0:192] cby_0__1__3_chany_bottom_out;
wire [0:192] cby_0__1__3_chany_top_out;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_0__2__0_ccff_tail;
wire [0:192] cby_0__2__0_chany_bottom_out;
wire [0:192] cby_0__2__0_chany_top_out;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_;
wire [0:0] cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_;
wire [0:0] cby_0__2__1_ccff_tail;
wire [0:192] cby_0__2__1_chany_bottom_out;
wire [0:192] cby_0__2__1_chany_top_out;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_0__2__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_;
wire [0:0] cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_;
wire [0:0] cby_1__1__0_ccff_tail;
wire [0:192] cby_1__1__0_chany_bottom_out;
wire [0:192] cby_1__1__0_chany_top_out;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__10_ccff_tail;
wire [0:192] cby_1__1__10_chany_bottom_out;
wire [0:192] cby_1__1__10_chany_top_out;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__11_ccff_tail;
wire [0:192] cby_1__1__11_chany_bottom_out;
wire [0:192] cby_1__1__11_chany_top_out;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__12_ccff_tail;
wire [0:192] cby_1__1__12_chany_bottom_out;
wire [0:192] cby_1__1__12_chany_top_out;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__13_ccff_tail;
wire [0:192] cby_1__1__13_chany_bottom_out;
wire [0:192] cby_1__1__13_chany_top_out;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__1_ccff_tail;
wire [0:192] cby_1__1__1_chany_bottom_out;
wire [0:192] cby_1__1__1_chany_top_out;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__2_ccff_tail;
wire [0:192] cby_1__1__2_chany_bottom_out;
wire [0:192] cby_1__1__2_chany_top_out;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__3_ccff_tail;
wire [0:192] cby_1__1__3_chany_bottom_out;
wire [0:192] cby_1__1__3_chany_top_out;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__4_ccff_tail;
wire [0:192] cby_1__1__4_chany_bottom_out;
wire [0:192] cby_1__1__4_chany_top_out;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__5_ccff_tail;
wire [0:192] cby_1__1__5_chany_bottom_out;
wire [0:192] cby_1__1__5_chany_top_out;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__6_ccff_tail;
wire [0:192] cby_1__1__6_chany_bottom_out;
wire [0:192] cby_1__1__6_chany_top_out;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__7_ccff_tail;
wire [0:192] cby_1__1__7_chany_bottom_out;
wire [0:192] cby_1__1__7_chany_top_out;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__8_ccff_tail;
wire [0:192] cby_1__1__8_chany_bottom_out;
wire [0:192] cby_1__1__8_chany_top_out;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__1__9_ccff_tail;
wire [0:192] cby_1__1__9_chany_bottom_out;
wire [0:192] cby_1__1__9_chany_top_out;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__0_ccff_tail;
wire [0:192] cby_1__2__0_chany_bottom_out;
wire [0:192] cby_1__2__0_chany_top_out;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_;
wire [0:0] cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_1__2__1_ccff_tail;
wire [0:192] cby_1__2__1_chany_bottom_out;
wire [0:192] cby_1__2__1_chany_top_out;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_;
wire [0:0] cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_;
wire [0:0] cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_;
wire [0:0] cby_3__2__0_ccff_tail;
wire [0:192] cby_3__2__0_chany_bottom_out;
wire [0:192] cby_3__2__0_chany_top_out;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_;
wire [0:0] cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_;
wire [0:0] cby_3__2__1_ccff_tail;
wire [0:192] cby_3__2__1_chany_bottom_out;
wire [0:192] cby_3__2__1_chany_top_out;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_;
wire [0:0] cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_;
wire [0:0] cby_4__1__0_ccff_tail;
wire [0:192] cby_4__1__0_chany_bottom_out;
wire [0:192] cby_4__1__0_chany_top_out;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_4__1__1_ccff_tail;
wire [0:192] cby_4__1__1_chany_bottom_out;
wire [0:192] cby_4__1__1_chany_top_out;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_4__1__2_ccff_tail;
wire [0:192] cby_4__1__2_chany_bottom_out;
wire [0:192] cby_4__1__2_chany_top_out;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_4__1__3_ccff_tail;
wire [0:192] cby_4__1__3_chany_bottom_out;
wire [0:192] cby_4__1__3_chany_top_out;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_;
wire [0:0] cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_4__2__0_ccff_tail;
wire [0:192] cby_4__2__0_chany_bottom_out;
wire [0:192] cby_4__2__0_chany_top_out;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_;
wire [0:0] cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] cby_4__2__1_ccff_tail;
wire [0:192] cby_4__2__1_chany_bottom_out;
wire [0:192] cby_4__2__1_chany_top_out;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_;
wire [0:0] cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_;
wire [0:0] cby_4__2__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_;
wire [0:0] grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_0_ccff_tail;
wire [0:0] grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_10_ccff_tail;
wire [0:0] grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_11_ccff_tail;
wire [0:0] grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_12_ccff_tail;
wire [0:0] grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_13_ccff_tail;
wire [0:0] grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_14_ccff_tail;
wire [0:0] grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_15_ccff_tail;
wire [0:0] grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_16_ccff_tail;
wire [0:0] grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_17_ccff_tail;
wire [0:0] grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_18_ccff_tail;
wire [0:0] grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_19_ccff_tail;
wire [0:0] grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_1_ccff_tail;
wire [0:0] grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_2_ccff_tail;
wire [0:0] grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_4_ccff_tail;
wire [0:0] grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_5_ccff_tail;
wire [0:0] grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_6_ccff_tail;
wire [0:0] grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_7_ccff_tail;
wire [0:0] grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_8_ccff_tail;
wire [0:0] grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_;
wire [0:0] grid_clb_9_ccff_tail;
wire [0:0] grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_;
wire [0:0] grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_;
wire [0:0] grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_;
wire [0:0] grid_io_bottom_0_ccff_tail;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_ccff_tail;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_ccff_tail;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_ccff_tail;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_0_ccff_tail;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_1_ccff_tail;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_2_ccff_tail;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_3_ccff_tail;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_4_ccff_tail;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_left_5_ccff_tail;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_0_ccff_tail;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_1_ccff_tail;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_2_ccff_tail;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_3_ccff_tail;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_4_ccff_tail;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_right_5_ccff_tail;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_0_ccff_tail;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_1_ccff_tail;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_2_ccff_tail;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
wire [0:0] grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
wire [0:0] grid_io_top_3_ccff_tail;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
wire [0:0] grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
wire [0:0] grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_error_0_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
wire [0:0] grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
wire [0:0] grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
wire [0:0] grid_router_1__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_1__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
wire [0:0] grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
wire [0:0] grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_error_0_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
wire [0:0] grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
wire [0:0] grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
wire [0:0] grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
wire [0:0] grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_error_0_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
wire [0:0] grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
wire [0:0] grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
wire [0:0] grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
wire [0:0] grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_error_0_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
wire [0:0] grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
wire [0:0] grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
wire [0:0] grid_router_4__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] grid_router_4__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_;
wire [0:0] sb_0__0__0_ccff_tail;
wire [0:192] sb_0__0__0_chanx_right_out;
wire [0:192] sb_0__0__0_chany_top_out;
wire [0:0] sb_0__1__0_ccff_tail;
wire [0:192] sb_0__1__0_chanx_right_out;
wire [0:192] sb_0__1__0_chany_bottom_out;
wire [0:192] sb_0__1__0_chany_top_out;
wire [0:0] sb_0__1__1_ccff_tail;
wire [0:192] sb_0__1__1_chanx_right_out;
wire [0:192] sb_0__1__1_chany_bottom_out;
wire [0:192] sb_0__1__1_chany_top_out;
wire [0:0] sb_0__2__0_ccff_tail;
wire [0:192] sb_0__2__0_chanx_right_out;
wire [0:192] sb_0__2__0_chany_bottom_out;
wire [0:192] sb_0__2__0_chany_top_out;
wire [0:0] sb_0__2__1_ccff_tail;
wire [0:192] sb_0__2__1_chanx_right_out;
wire [0:192] sb_0__2__1_chany_bottom_out;
wire [0:192] sb_0__2__1_chany_top_out;
wire [0:0] sb_0__3__0_ccff_tail;
wire [0:192] sb_0__3__0_chanx_right_out;
wire [0:192] sb_0__3__0_chany_bottom_out;
wire [0:192] sb_0__3__0_chany_top_out;
wire [0:0] sb_0__6__0_ccff_tail;
wire [0:192] sb_0__6__0_chanx_right_out;
wire [0:192] sb_0__6__0_chany_bottom_out;
wire [0:0] sb_1__0__0_ccff_tail;
wire [0:192] sb_1__0__0_chanx_left_out;
wire [0:192] sb_1__0__0_chanx_right_out;
wire [0:192] sb_1__0__0_chany_top_out;
wire [0:0] sb_1__0__1_ccff_tail;
wire [0:192] sb_1__0__1_chanx_left_out;
wire [0:192] sb_1__0__1_chanx_right_out;
wire [0:192] sb_1__0__1_chany_top_out;
wire [0:0] sb_1__0__2_ccff_tail;
wire [0:192] sb_1__0__2_chanx_left_out;
wire [0:192] sb_1__0__2_chanx_right_out;
wire [0:192] sb_1__0__2_chany_top_out;
wire [0:0] sb_1__1__0_ccff_tail;
wire [0:192] sb_1__1__0_chanx_left_out;
wire [0:192] sb_1__1__0_chanx_right_out;
wire [0:192] sb_1__1__0_chany_bottom_out;
wire [0:192] sb_1__1__0_chany_top_out;
wire [0:0] sb_1__1__1_ccff_tail;
wire [0:192] sb_1__1__1_chanx_left_out;
wire [0:192] sb_1__1__1_chanx_right_out;
wire [0:192] sb_1__1__1_chany_bottom_out;
wire [0:192] sb_1__1__1_chany_top_out;
wire [0:0] sb_1__2__0_ccff_tail;
wire [0:192] sb_1__2__0_chanx_left_out;
wire [0:192] sb_1__2__0_chanx_right_out;
wire [0:192] sb_1__2__0_chany_bottom_out;
wire [0:192] sb_1__2__0_chany_top_out;
wire [0:0] sb_1__2__1_ccff_tail;
wire [0:192] sb_1__2__1_chanx_left_out;
wire [0:192] sb_1__2__1_chanx_right_out;
wire [0:192] sb_1__2__1_chany_bottom_out;
wire [0:192] sb_1__2__1_chany_top_out;
wire [0:0] sb_1__3__0_ccff_tail;
wire [0:192] sb_1__3__0_chanx_left_out;
wire [0:192] sb_1__3__0_chanx_right_out;
wire [0:192] sb_1__3__0_chany_bottom_out;
wire [0:192] sb_1__3__0_chany_top_out;
wire [0:0] sb_1__3__1_ccff_tail;
wire [0:192] sb_1__3__1_chanx_left_out;
wire [0:192] sb_1__3__1_chanx_right_out;
wire [0:192] sb_1__3__1_chany_bottom_out;
wire [0:192] sb_1__3__1_chany_top_out;
wire [0:0] sb_1__3__2_ccff_tail;
wire [0:192] sb_1__3__2_chanx_left_out;
wire [0:192] sb_1__3__2_chanx_right_out;
wire [0:192] sb_1__3__2_chany_bottom_out;
wire [0:192] sb_1__3__2_chany_top_out;
wire [0:0] sb_1__3__3_ccff_tail;
wire [0:192] sb_1__3__3_chanx_left_out;
wire [0:192] sb_1__3__3_chanx_right_out;
wire [0:192] sb_1__3__3_chany_bottom_out;
wire [0:192] sb_1__3__3_chany_top_out;
wire [0:0] sb_1__3__4_ccff_tail;
wire [0:192] sb_1__3__4_chanx_left_out;
wire [0:192] sb_1__3__4_chanx_right_out;
wire [0:192] sb_1__3__4_chany_bottom_out;
wire [0:192] sb_1__3__4_chany_top_out;
wire [0:0] sb_1__3__5_ccff_tail;
wire [0:192] sb_1__3__5_chanx_left_out;
wire [0:192] sb_1__3__5_chanx_right_out;
wire [0:192] sb_1__3__5_chany_bottom_out;
wire [0:192] sb_1__3__5_chany_top_out;
wire [0:0] sb_1__3__6_ccff_tail;
wire [0:192] sb_1__3__6_chanx_left_out;
wire [0:192] sb_1__3__6_chanx_right_out;
wire [0:192] sb_1__3__6_chany_bottom_out;
wire [0:192] sb_1__3__6_chany_top_out;
wire [0:0] sb_1__6__0_ccff_tail;
wire [0:192] sb_1__6__0_chanx_left_out;
wire [0:192] sb_1__6__0_chanx_right_out;
wire [0:192] sb_1__6__0_chany_bottom_out;
wire [0:0] sb_1__6__1_ccff_tail;
wire [0:192] sb_1__6__1_chanx_left_out;
wire [0:192] sb_1__6__1_chanx_right_out;
wire [0:192] sb_1__6__1_chany_bottom_out;
wire [0:0] sb_1__6__2_ccff_tail;
wire [0:192] sb_1__6__2_chanx_left_out;
wire [0:192] sb_1__6__2_chanx_right_out;
wire [0:192] sb_1__6__2_chany_bottom_out;
wire [0:0] sb_3__1__0_ccff_tail;
wire [0:192] sb_3__1__0_chanx_left_out;
wire [0:192] sb_3__1__0_chanx_right_out;
wire [0:192] sb_3__1__0_chany_bottom_out;
wire [0:192] sb_3__1__0_chany_top_out;
wire [0:0] sb_3__1__1_ccff_tail;
wire [0:192] sb_3__1__1_chanx_left_out;
wire [0:192] sb_3__1__1_chanx_right_out;
wire [0:192] sb_3__1__1_chany_bottom_out;
wire [0:192] sb_3__1__1_chany_top_out;
wire [0:0] sb_3__2__0_ccff_tail;
wire [0:192] sb_3__2__0_chanx_left_out;
wire [0:192] sb_3__2__0_chanx_right_out;
wire [0:192] sb_3__2__0_chany_bottom_out;
wire [0:192] sb_3__2__0_chany_top_out;
wire [0:0] sb_3__2__1_ccff_tail;
wire [0:192] sb_3__2__1_chanx_left_out;
wire [0:192] sb_3__2__1_chanx_right_out;
wire [0:192] sb_3__2__1_chany_bottom_out;
wire [0:192] sb_3__2__1_chany_top_out;
wire [0:0] sb_4__0__0_ccff_tail;
wire [0:192] sb_4__0__0_chanx_left_out;
wire [0:192] sb_4__0__0_chany_top_out;
wire [0:0] sb_4__1__0_ccff_tail;
wire [0:192] sb_4__1__0_chanx_left_out;
wire [0:192] sb_4__1__0_chany_bottom_out;
wire [0:192] sb_4__1__0_chany_top_out;
wire [0:0] sb_4__1__1_ccff_tail;
wire [0:192] sb_4__1__1_chanx_left_out;
wire [0:192] sb_4__1__1_chany_bottom_out;
wire [0:192] sb_4__1__1_chany_top_out;
wire [0:0] sb_4__2__0_ccff_tail;
wire [0:192] sb_4__2__0_chanx_left_out;
wire [0:192] sb_4__2__0_chany_bottom_out;
wire [0:192] sb_4__2__0_chany_top_out;
wire [0:0] sb_4__2__1_ccff_tail;
wire [0:192] sb_4__2__1_chanx_left_out;
wire [0:192] sb_4__2__1_chany_bottom_out;
wire [0:192] sb_4__2__1_chany_top_out;
wire [0:0] sb_4__3__0_ccff_tail;
wire [0:192] sb_4__3__0_chanx_left_out;
wire [0:192] sb_4__3__0_chany_bottom_out;
wire [0:192] sb_4__3__0_chany_top_out;
wire [0:0] sb_4__6__0_ccff_tail;
wire [0:192] sb_4__6__0_chanx_left_out;
wire [0:192] sb_4__6__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top grid_io_top_1__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__6__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__6__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__6__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_4__7_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__6__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_right grid_io_right_5__6_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_5__5_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_5__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_5__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_right grid_io_right_5__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_4_ccff_tail));

	grid_io_right grid_io_right_5__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_5_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__2__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[128:135]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[136:143]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	grid_io_left grid_io_left_0__5_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[144:151]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__2__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_4_ccff_tail));

	grid_io_left grid_io_left_0__6_ (
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[152:159]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_5_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_2__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_3__2__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__5__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_3__2__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_1__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_4__1_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_4__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_4__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_4__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_4__6_ (
		.prog_clk(prog_clk),
		.set(set),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__6__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.ccff_head(cby_4__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_router grid_router_1__2_ (
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_router_1__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_0_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_4_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.left_width_0_height_0_subtile_0__pin_router_address_2_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.right_width_0_height_0_subtile_0__pin_error_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_error_0_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_));

	grid_router grid_router_1__5_ (
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_router_1__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_0_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_4_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.left_width_0_height_0_subtile_0__pin_router_address_2_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.right_width_0_height_0_subtile_0__pin_error_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_error_0_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_));

	grid_router grid_router_4__2_ (
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_router_4__2__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.left_width_0_height_0_subtile_0__pin_router_address_2_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.right_width_0_height_0_subtile_0__pin_error_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_error_0_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_));

	grid_router grid_router_4__5_ (
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.top_width_0_height_0_subtile_0__pin_clk_0_(grid_router_4__5__undriven_top_width_0_height_0_subtile_0__pin_clk_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.right_width_0_height_0_subtile_0__pin_router_address_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.left_width_0_height_0_subtile_0__pin_router_address_2_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.right_width_0_height_0_subtile_0__pin_error_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_error_0_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_));

	sb_0__0_ sb_0__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:192]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:192]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__2__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:192]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__2__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_5_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:192]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__2_ sb_0__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__0_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.chany_bottom_in(cby_0__2__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_0_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_0_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__2__0_chany_top_out[0:192]),
		.chanx_right_out(sb_0__2__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__2__0_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__2__0_ccff_tail));

	sb_0__2_ sb_0__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__1_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.chany_bottom_in(cby_0__2__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_1_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_1_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_4_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__6__0_ccff_tail),
		.chany_top_out(sb_0__2__1_chany_top_out[0:192]),
		.chanx_right_out(sb_0__2__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__2__1_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__2__1_ccff_tail));

	sb_0__3_ sb_0__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__0_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_4_ccff_tail),
		.chany_top_out(sb_0__3__0_chany_top_out[0:192]),
		.chanx_right_out(sb_0__3__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__3__0_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__3__0_ccff_tail));

	sb_0__6_ sb_0__6_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__0_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_5_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__6__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_0__6__0_chany_bottom_out[0:192]),
		.ccff_tail(sb_0__6__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:192]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:192]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:192]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:192]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:192]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:192]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:192]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:192]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:192]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_error_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__1_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_0_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:192]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:192]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__2__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_error_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__4_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_1_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:192]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:192]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__2_ sb_1__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__2_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__2__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_0_right_width_0_height_0_subtile_0__pin_error_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_0_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_0_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.chanx_left_in(cbx_1__2__0_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_0_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_0_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.ccff_head(cby_1__2__0_ccff_tail),
		.chany_top_out(sb_1__2__0_chany_top_out[0:192]),
		.chanx_right_out(sb_1__2__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__2__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__2__0_chanx_left_out[0:192]),
		.ccff_tail(sb_1__2__0_ccff_tail));

	sb_1__2_ sb_1__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__5_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__2__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_1_right_width_0_height_0_subtile_0__pin_error_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_1_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_1_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.chanx_left_in(cbx_1__2__1_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_1_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_1_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__2__1_chany_top_out[0:192]),
		.chanx_right_out(sb_1__2__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__2__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__2__1_chanx_left_out[0:192]),
		.ccff_tail(sb_1__2__1_ccff_tail));

	sb_1__3_ sb_1__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__3_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__0_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__3__0_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__0_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__0_ccff_tail));

	sb_1__3_ sb_2__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__6_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__1_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__3__1_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__1_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__1_ccff_tail));

	sb_1__3_ sb_2__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__7_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__2_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__3__2_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__2_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__2_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__2_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__2_ccff_tail));

	sb_1__3_ sb_2__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__8_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__3_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__3__3_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__3_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__3_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__3_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__3_ccff_tail));

	sb_1__3_ sb_2__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__9_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__4_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(cby_1__2__1_ccff_tail),
		.chany_top_out(sb_1__3__4_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__4_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__4_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__4_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__4_ccff_tail));

	sb_1__3_ sb_2__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__10_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__5_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__3__5_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__5_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__5_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__5_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__5_ccff_tail));

	sb_1__3_ sb_3__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__3__11_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__8_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__3__6_chany_top_out[0:192]),
		.chanx_right_out(sb_1__3__6_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__3__6_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__3__6_chanx_left_out[0:192]),
		.ccff_tail(sb_1__3__6_ccff_tail));

	sb_1__6_ sb_1__6_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__1_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__6__0_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__6__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__6__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__6__0_chanx_left_out[0:192]),
		.ccff_tail(sb_1__6__0_ccff_tail));

	sb_1__6_ sb_2__6_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__2_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__6__1_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__6__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__6__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__6__1_chanx_left_out[0:192]),
		.ccff_tail(sb_1__6__1_ccff_tail));

	sb_1__6_ sb_3__6_ (
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__6__3_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__6__2_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chanx_right_out(sb_1__6__2_chanx_right_out[0:192]),
		.chany_bottom_out(sb_1__6__2_chany_bottom_out[0:192]),
		.chanx_left_out(sb_1__6__2_chanx_left_out[0:192]),
		.ccff_tail(sb_1__6__2_ccff_tail));

	sb_3__1_ sb_3__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__6_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(cby_4__2__0_ccff_tail),
		.chany_top_out(sb_3__1__0_chany_top_out[0:192]),
		.chanx_right_out(sb_3__1__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_3__1__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_3__1__0_chanx_left_out[0:192]),
		.ccff_tail(sb_3__1__0_ccff_tail));

	sb_3__1_ sb_3__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_3__2__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_left_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__9_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_3__1__1_chany_top_out[0:192]),
		.chanx_right_out(sb_3__1__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_3__1__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_3__1__1_chanx_left_out[0:192]),
		.ccff_tail(sb_3__1__1_ccff_tail));

	sb_3__2_ sb_3__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__2_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.chany_bottom_in(cby_3__2__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_2_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_2_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__7_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_3__2__0_chany_top_out[0:192]),
		.chanx_right_out(sb_3__2__0_chanx_right_out[0:192]),
		.chany_bottom_out(sb_3__2__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_3__2__0_chanx_left_out[0:192]),
		.ccff_tail(sb_3__2__0_ccff_tail));

	sb_3__2_ sb_3__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_left_width_0_height_0_subtile_0__pin_O_1_),
		.chanx_right_in(cbx_1__2__3_chanx_left_out[0:192]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.chany_bottom_in(cby_3__2__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_9_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_13_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_17_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_21_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_25_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_29_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_33_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_37_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_41_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_45_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_49_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_53_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_57_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_61_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_65_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_69_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_73_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_77_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_81_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_85_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_89_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_93_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_97_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_101_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_105_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_109_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_113_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_117_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_121_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_125_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_129_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_133_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_137_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_141_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_145_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_149_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_153_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_157_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_161_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_165_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_169_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_173_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_177_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_181_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_185_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_189_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_193_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_197_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_201_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_205_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_209_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_213_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_217_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_221_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_225_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_229_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_233_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_237_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_241_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_245_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_249_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_253_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_257_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_261_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_265_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_269_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_273_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_277_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_281_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_285_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_289_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_293_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_297_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_301_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_305_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_309_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_313_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_317_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_321_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_325_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_329_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_333_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_(grid_router_3_left_width_0_height_0_subtile_0__pin_channel_out_op_337_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_(grid_router_3_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__10_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_3__2__1_chany_top_out[0:192]),
		.chanx_right_out(sb_3__2__1_chanx_right_out[0:192]),
		.chany_bottom_out(sb_3__2__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_3__2__1_chanx_left_out[0:192]),
		.ccff_tail(sb_3__2__1_ccff_tail));

	sb_4__0_ sb_4__0_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_4__0__0_chany_top_out[0:192]),
		.chanx_left_out(sb_4__0__0_chanx_left_out[0:192]),
		.ccff_tail(sb_4__0__0_ccff_tail));

	sb_4__1_ sb_4__1_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__2__0_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_error_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_5_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_2_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_4__1__0_chany_top_out[0:192]),
		.chany_bottom_out(sb_4__1__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__1__0_chanx_left_out[0:192]),
		.ccff_tail(sb_4__1__0_ccff_tail));

	sb_4__1_ sb_4__4_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__2__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_error_0_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__2_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_(grid_router_3_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_4__1__1_chany_top_out[0:192]),
		.chany_bottom_out(sb_4__1__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__1__1_chanx_left_out[0:192]),
		.ccff_tail(sb_4__1__1_ccff_tail));

	sb_4__2_ sb_4__2_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__1_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__2__0_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_4_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_2_right_width_0_height_0_subtile_0__pin_error_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_2_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_2_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.chanx_left_in(cbx_1__2__2_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_2_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_2_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_4__2__0_chany_top_out[0:192]),
		.chany_bottom_out(sb_4__2__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__2__0_chanx_left_out[0:192]),
		.ccff_tail(sb_4__2__0_ccff_tail));

	sb_4__2_ sb_4__5_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__3_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__2__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_(grid_router_3_right_width_0_height_0_subtile_0__pin_error_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_15_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_19_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_23_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_27_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_31_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_35_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_39_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_43_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_47_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_51_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_55_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_59_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_63_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_67_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_71_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_75_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_79_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_83_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_87_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_91_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_95_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_99_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_103_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_107_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_111_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_115_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_119_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_123_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_127_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_131_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_135_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_139_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_143_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_147_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_151_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_155_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_159_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_163_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_167_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_171_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_175_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_179_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_183_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_187_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_191_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_195_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_199_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_203_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_207_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_211_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_215_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_219_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_223_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_227_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_231_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_235_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_239_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_243_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_247_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_251_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_255_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_259_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_263_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_267_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_271_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_275_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_279_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_283_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_287_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_291_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_295_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_299_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_303_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_307_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_311_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_315_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_319_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_323_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_327_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_331_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_335_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_(grid_router_3_right_width_0_height_0_subtile_0__pin_channel_out_op_339_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_(grid_router_3_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_),
		.chanx_left_in(cbx_1__2__3_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_10_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_14_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_18_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_22_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_26_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_30_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_34_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_38_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_42_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_46_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_50_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_54_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_58_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_62_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_66_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_70_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_74_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_78_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_82_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_86_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_90_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_94_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_98_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_102_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_106_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_110_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_114_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_118_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_122_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_126_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_130_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_134_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_138_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_142_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_146_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_150_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_154_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_158_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_162_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_166_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_170_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_174_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_178_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_182_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_186_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_190_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_194_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_198_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_202_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_206_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_210_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_214_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_218_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_222_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_226_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_230_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_234_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_238_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_242_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_246_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_250_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_254_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_258_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_262_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_266_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_270_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_274_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_278_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_282_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_286_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_290_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_294_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_298_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_302_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_306_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_310_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_314_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_318_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_322_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_326_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_330_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_334_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_(grid_router_3_top_width_0_height_0_subtile_0__pin_channel_out_op_338_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_(grid_router_3_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_),
		.ccff_head(cby_4__2__1_ccff_tail),
		.chany_top_out(sb_4__2__1_chany_top_out[0:192]),
		.chany_bottom_out(sb_4__2__1_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__2__1_chanx_left_out[0:192]),
		.ccff_tail(sb_4__2__1_ccff_tail));

	sb_4__3_ sb_4__3_ (
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__2_chany_bottom_out[0:192]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__1_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__3__11_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_4__3__0_chany_top_out[0:192]),
		.chany_bottom_out(sb_4__3__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__3__0_chanx_left_out[0:192]),
		.ccff_tail(sb_4__3__0_ccff_tail));

	sb_4__6_ sb_4__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__1__3_chany_top_out[0:192]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_3_),
		.chanx_left_in(cbx_1__6__3_chanx_right_out[0:192]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_4__6__0_chany_bottom_out[0:192]),
		.chanx_left_out(sb_4__6__0_chanx_left_out[0:192]),
		.ccff_tail(sb_4__6__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:192]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:192]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:192]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__0__0_chanx_left_out[0:192]),
		.ccff_head(sb_4__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:192]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:192]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__1__0_chanx_left_out[0:192]),
		.ccff_head(sb_4__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_4__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__1__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__1__1_chanx_left_out[0:192]),
		.ccff_head(sb_4__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_1_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_router_address_5_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_7_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_11_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_15_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_19_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_23_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_27_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_31_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_35_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_39_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_43_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_47_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_51_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_55_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_59_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_63_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_67_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_71_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_75_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_79_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_83_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_87_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_91_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_95_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_99_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_103_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_107_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_111_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_115_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_119_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_123_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_127_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_131_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_135_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_139_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_143_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_147_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_151_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_155_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_159_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_163_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_167_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_171_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_175_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_179_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_183_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_187_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_191_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_195_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_199_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_203_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_207_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_211_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_215_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_219_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_223_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_227_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_231_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_235_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_239_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_243_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_247_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_251_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_255_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_259_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_263_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_267_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_271_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_275_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_279_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_283_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_287_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_291_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_295_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_299_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_303_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_307_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_311_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_315_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_319_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_323_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_327_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_331_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_335_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_in_ip_339_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_3_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_7_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__2_ cbx_1__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__2__0_chanx_left_out[0:192]),
		.ccff_head(sb_1__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__0_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__2__0_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__0_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.ccff_tail(cbx_1__2__0_ccff_tail));

	cbx_1__2_ cbx_1__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__2__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__2__1_chanx_left_out[0:192]),
		.ccff_head(sb_1__2__1_ccff_tail),
		.chanx_left_out(cbx_1__2__1_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__2__1_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__1_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.ccff_tail(cbx_1__2__1_ccff_tail));

	cbx_1__2_ cbx_4__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__2__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__2__0_chanx_left_out[0:192]),
		.ccff_head(sb_4__2__0_ccff_tail),
		.chanx_left_out(cbx_1__2__2_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__2__2_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__2_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.ccff_tail(cbx_1__2__2_ccff_tail));

	cbx_1__2_ cbx_4__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_3__2__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__2__1_chanx_left_out[0:192]),
		.ccff_head(sb_4__2__1_ccff_tail),
		.chanx_left_out(cbx_1__2__3_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__2__3_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__2__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_reset_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_router_address_3_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_9_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_13_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_17_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_21_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_25_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_29_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_33_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_37_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_41_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_45_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_49_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_53_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_57_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_61_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_65_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_69_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_73_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_77_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_81_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_85_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_89_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_93_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_97_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_101_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_105_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_109_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_113_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_117_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_121_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_125_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_129_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_133_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_137_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_141_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_145_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_149_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_153_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_157_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_161_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_165_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_169_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_173_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_177_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_181_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_185_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_189_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_193_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_197_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_201_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_205_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_209_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_213_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_217_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_221_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_225_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_229_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_233_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_237_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_241_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_245_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_249_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_253_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_257_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_261_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_265_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_269_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_273_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_277_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_281_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_285_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_289_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_293_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_297_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_301_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_305_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_309_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_313_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_317_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_321_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_325_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_329_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_333_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_in_ip_337_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_5_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_(cbx_1__2__3_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_9_),
		.ccff_tail(cbx_1__2__3_ccff_tail));

	cbx_1__3_ cbx_1__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__3__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__0_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__0_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__0_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__0_ccff_tail));

	cbx_1__3_ cbx_2__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__1_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__1_ccff_tail),
		.chanx_left_out(cbx_1__3__1_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__1_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__1_ccff_tail));

	cbx_1__3_ cbx_2__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__2_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__2_ccff_tail),
		.chanx_left_out(cbx_1__3__2_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__2_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__2_ccff_tail));

	cbx_1__3_ cbx_2__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__3_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__3_ccff_tail),
		.chanx_left_out(cbx_1__3__3_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__3_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__3_ccff_tail));

	cbx_1__3_ cbx_2__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__4_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__4_ccff_tail),
		.chanx_left_out(cbx_1__3__4_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__4_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__4_ccff_tail));

	cbx_1__3_ cbx_2__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__2__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__5_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__5_ccff_tail),
		.chanx_left_out(cbx_1__3__5_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__5_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__5_ccff_tail));

	cbx_1__3_ cbx_3__1_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_3__1__0_chanx_left_out[0:192]),
		.ccff_head(sb_3__1__0_ccff_tail),
		.chanx_left_out(cbx_1__3__6_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__6_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__6_ccff_tail));

	cbx_1__3_ cbx_3__2_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__2_chanx_right_out[0:192]),
		.chanx_right_in(sb_3__2__0_chanx_left_out[0:192]),
		.ccff_head(sb_3__2__0_ccff_tail),
		.chanx_left_out(cbx_1__3__7_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__7_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__7_ccff_tail));

	cbx_1__3_ cbx_3__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__3_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__3__6_chanx_left_out[0:192]),
		.ccff_head(sb_1__3__6_ccff_tail),
		.chanx_left_out(cbx_1__3__8_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__8_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__8_ccff_tail));

	cbx_1__3_ cbx_3__4_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__4_chanx_right_out[0:192]),
		.chanx_right_in(sb_3__1__1_chanx_left_out[0:192]),
		.ccff_head(sb_3__1__1_ccff_tail),
		.chanx_left_out(cbx_1__3__9_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__9_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__9_ccff_tail));

	cbx_1__3_ cbx_3__5_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__5_chanx_right_out[0:192]),
		.chanx_right_in(sb_3__2__1_chanx_left_out[0:192]),
		.ccff_head(sb_3__2__1_ccff_tail),
		.chanx_left_out(cbx_1__3__10_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__10_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__10_ccff_tail));

	cbx_1__3_ cbx_4__3_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__3__6_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__3__0_chanx_left_out[0:192]),
		.ccff_head(sb_4__3__0_ccff_tail),
		.chanx_left_out(cbx_1__3__11_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__3__11_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__3__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__3__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__3__11_ccff_tail));

	cbx_1__6_ cbx_1__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__6__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__6__0_chanx_left_out[0:192]),
		.ccff_head(sb_1__6__0_ccff_tail),
		.chanx_left_out(cbx_1__6__0_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__6__0_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__6__0_ccff_tail));

	cbx_1__6_ cbx_2__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__6__0_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__6__1_chanx_left_out[0:192]),
		.ccff_head(sb_1__6__1_ccff_tail),
		.chanx_left_out(cbx_1__6__1_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__6__1_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__6__1_ccff_tail));

	cbx_1__6_ cbx_3__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__6__1_chanx_right_out[0:192]),
		.chanx_right_in(sb_1__6__2_chanx_left_out[0:192]),
		.ccff_head(sb_1__6__2_ccff_tail),
		.chanx_left_out(cbx_1__6__2_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__6__2_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__6__2_ccff_tail));

	cbx_1__6_ cbx_4__6_ (
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__6__2_chanx_right_out[0:192]),
		.chanx_right_in(sb_4__6__0_chanx_left_out[0:192]),
		.ccff_head(sb_4__6__0_ccff_tail),
		.chanx_left_out(cbx_1__6__3_chanx_left_out[0:192]),
		.chanx_right_out(cbx_1__6__3_chanx_right_out[0:192]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__6__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__6__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.ccff_tail(cbx_1__6__3_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:192]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:192]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__2__0_chany_top_out[0:192]),
		.chany_top_in(sb_0__3__0_chany_bottom_out[0:192]),
		.ccff_head(sb_0__2__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__3__0_chany_top_out[0:192]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:192]),
		.ccff_head(sb_0__3__0_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__2__1_chany_top_out[0:192]),
		.chany_top_in(sb_0__6__0_chany_bottom_out[0:192]),
		.ccff_head(sb_0__2__1_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__2_ cby_0__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:192]),
		.chany_top_in(sb_0__2__0_chany_bottom_out[0:192]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__2__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__2__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_0__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__2__0_ccff_tail));

	cby_0__2_ cby_0__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:192]),
		.chany_top_in(sb_0__2__1_chany_bottom_out[0:192]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__2__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_0__2__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_0__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__2__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__2__1_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:192]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__0_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__2__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__0_chany_top_out[0:192]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__0_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__2__1_chany_top_out[0:192]),
		.chany_top_in(sb_1__6__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__2__1_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__1_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__2_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__1_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__2_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__3_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__2_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_2__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__3_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__4_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__3_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_2__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__4_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__5_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__4_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_2__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__5_chany_top_out[0:192]),
		.chany_top_in(sb_1__6__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__5_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_3__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:192]),
		.chany_top_in(sb_3__1__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_3__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__0_chany_top_out[0:192]),
		.chany_top_in(sb_1__3__6_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__7_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_1__1_ cby_3__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__3__6_chany_top_out[0:192]),
		.chany_top_in(sb_3__1__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__8_ccff_tail),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__12_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__12_ccff_tail));

	cby_1__1_ cby_3__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__2__1_chany_top_out[0:192]),
		.chany_top_in(sb_1__6__2_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__10_ccff_tail),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__13_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_1__1__13_ccff_tail));

	cby_1__2_ cby_1__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:192]),
		.chany_top_in(sb_1__2__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__2__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__2__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_1__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.ccff_tail(cby_1__2__0_ccff_tail));

	cby_1__2_ cby_1__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:192]),
		.chany_top_in(sb_1__2__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__2__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_1__2__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__2__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_1__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.ccff_tail(cby_1__2__1_ccff_tail));

	cby_3__2_ cby_3__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__0_chany_top_out[0:192]),
		.chany_top_in(sb_3__2__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__6_ccff_tail),
		.chany_bottom_out(cby_3__2__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_3__2__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_3__2__0_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_3__2__0_ccff_tail));

	cby_3__2_ cby_3__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_3__1__1_chany_top_out[0:192]),
		.chany_top_in(sb_3__2__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__9_ccff_tail),
		.chany_bottom_out(cby_3__2__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_3__2__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_router_address_2_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_8_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_12_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_16_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_20_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_24_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_28_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_32_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_36_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_40_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_44_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_48_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_52_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_56_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_60_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_64_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_68_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_72_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_76_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_80_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_84_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_88_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_92_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_96_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_100_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_104_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_108_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_112_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_116_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_120_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_124_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_128_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_132_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_136_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_140_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_144_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_148_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_152_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_156_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_160_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_164_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_168_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_172_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_176_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_180_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_184_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_188_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_192_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_196_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_200_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_204_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_208_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_212_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_216_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_220_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_224_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_228_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_232_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_236_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_240_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_244_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_248_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_252_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_256_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_260_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_264_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_268_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_272_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_276_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_280_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_284_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_288_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_292_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_296_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_300_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_304_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_308_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_312_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_316_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_320_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_324_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_328_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_332_),
		.right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_channel_in_ip_336_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_0_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_4_),
		.right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_(cby_3__2__1_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_8_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_3__2__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_3__2__1_ccff_tail));

	cby_4__1_ cby_4__1_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__0__0_chany_top_out[0:192]),
		.chany_top_in(sb_4__1__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_4__1__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__1__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_4__1__0_ccff_tail));

	cby_4__1_ cby_4__3_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__2__0_chany_top_out[0:192]),
		.chany_top_in(sb_4__3__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__2__2_ccff_tail),
		.chany_bottom_out(cby_4__1__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__1__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_4__1__1_ccff_tail));

	cby_4__1_ cby_4__4_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__3__0_chany_top_out[0:192]),
		.chany_top_in(sb_4__1__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__3__11_ccff_tail),
		.chany_bottom_out(cby_4__1__2_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__1__2_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_4__1__2_ccff_tail));

	cby_4__1_ cby_4__6_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__2__1_chany_top_out[0:192]),
		.chany_top_in(sb_4__6__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__2__3_ccff_tail),
		.chany_bottom_out(cby_4__1__3_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__1__3_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.ccff_tail(cby_4__1__3_ccff_tail));

	cby_4__2_ cby_4__2_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__0_chany_top_out[0:192]),
		.chany_top_in(sb_4__2__0_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_4__2__0_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__2__0_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__2__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_4__2__0_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.ccff_tail(cby_4__2__0_ccff_tail));

	cby_4__2_ cby_4__5_ (
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__1_chany_top_out[0:192]),
		.chany_top_in(sb_4__2__1_chany_bottom_out[0:192]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_4__2__1_chany_bottom_out[0:192]),
		.chany_top_out(cby_4__2__1_chany_top_out[0:192]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__2__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_router_address_4_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_6_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_10_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_14_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_18_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_22_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_26_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_30_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_34_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_38_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_42_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_46_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_50_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_54_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_58_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_62_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_66_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_70_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_74_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_78_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_82_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_86_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_90_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_94_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_98_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_102_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_106_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_110_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_114_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_118_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_122_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_126_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_130_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_134_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_138_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_142_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_146_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_150_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_154_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_158_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_162_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_166_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_170_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_174_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_178_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_182_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_186_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_190_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_194_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_198_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_202_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_206_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_210_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_214_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_218_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_222_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_226_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_230_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_234_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_238_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_242_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_246_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_250_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_254_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_258_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_262_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_266_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_270_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_274_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_278_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_282_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_286_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_290_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_294_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_298_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_302_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_306_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_310_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_314_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_318_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_322_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_326_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_330_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_334_),
		.left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_channel_in_ip_338_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_2_),
		.left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_(cby_4__2__1_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_in_op_6_),
		.ccff_tail(cby_4__2__1_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype wire




