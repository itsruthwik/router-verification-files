//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jun 28 12:51:27 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__1_ -----
module sb_0__1_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:192] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
//----- INPUT PORTS -----
input [0:192] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:192] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:192] chany_top_out;
//----- OUTPUT PORTS -----
output [0:192] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:192] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_10_sram;
wire [0:3] mux_tree_tapbuf_size10_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_11_sram;
wire [0:3] mux_tree_tapbuf_size10_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_12_sram;
wire [0:3] mux_tree_tapbuf_size10_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_13_sram;
wire [0:3] mux_tree_tapbuf_size10_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_14_sram;
wire [0:3] mux_tree_tapbuf_size10_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_15_sram;
wire [0:3] mux_tree_tapbuf_size10_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_1_sram;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_2_sram;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_3_sram;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_4_sram;
wire [0:3] mux_tree_tapbuf_size10_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_5_sram;
wire [0:3] mux_tree_tapbuf_size10_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_6_sram;
wire [0:3] mux_tree_tapbuf_size10_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_7_sram;
wire [0:3] mux_tree_tapbuf_size10_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_8_sram;
wire [0:3] mux_tree_tapbuf_size10_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_9_sram;
wire [0:3] mux_tree_tapbuf_size10_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_11_sram;
wire [0:3] mux_tree_tapbuf_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_12_sram;
wire [0:3] mux_tree_tapbuf_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_13_sram;
wire [0:3] mux_tree_tapbuf_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_14_sram;
wire [0:3] mux_tree_tapbuf_size11_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_15_sram;
wire [0:3] mux_tree_tapbuf_size11_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_16_sram;
wire [0:3] mux_tree_tapbuf_size11_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_17_sram;
wire [0:3] mux_tree_tapbuf_size11_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_18_sram;
wire [0:3] mux_tree_tapbuf_size11_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_19_sram;
wire [0:3] mux_tree_tapbuf_size11_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_20_sram;
wire [0:3] mux_tree_tapbuf_size11_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_21_sram;
wire [0:3] mux_tree_tapbuf_size11_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_22_sram;
wire [0:3] mux_tree_tapbuf_size11_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_23_sram;
wire [0:3] mux_tree_tapbuf_size11_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_24_sram;
wire [0:3] mux_tree_tapbuf_size11_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_25_sram;
wire [0:3] mux_tree_tapbuf_size11_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_26_sram;
wire [0:3] mux_tree_tapbuf_size11_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_27_sram;
wire [0:3] mux_tree_tapbuf_size11_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_28_sram;
wire [0:3] mux_tree_tapbuf_size11_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_29_sram;
wire [0:3] mux_tree_tapbuf_size11_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_30_sram;
wire [0:3] mux_tree_tapbuf_size11_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_31_sram;
wire [0:3] mux_tree_tapbuf_size11_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_32_sram;
wire [0:3] mux_tree_tapbuf_size11_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_33_sram;
wire [0:3] mux_tree_tapbuf_size11_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_34_sram;
wire [0:3] mux_tree_tapbuf_size11_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_35_sram;
wire [0:3] mux_tree_tapbuf_size11_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_36_sram;
wire [0:3] mux_tree_tapbuf_size11_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_37_sram;
wire [0:3] mux_tree_tapbuf_size11_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_38_sram;
wire [0:3] mux_tree_tapbuf_size11_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_39_sram;
wire [0:3] mux_tree_tapbuf_size11_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_40_sram;
wire [0:3] mux_tree_tapbuf_size11_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_41_sram;
wire [0:3] mux_tree_tapbuf_size11_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_42_sram;
wire [0:3] mux_tree_tapbuf_size11_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_43_sram;
wire [0:3] mux_tree_tapbuf_size11_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_44_sram;
wire [0:3] mux_tree_tapbuf_size11_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_45_sram;
wire [0:3] mux_tree_tapbuf_size11_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_46_sram;
wire [0:3] mux_tree_tapbuf_size11_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_47_sram;
wire [0:3] mux_tree_tapbuf_size11_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_48_sram;
wire [0:3] mux_tree_tapbuf_size11_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_49_sram;
wire [0:3] mux_tree_tapbuf_size11_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_50_sram;
wire [0:3] mux_tree_tapbuf_size11_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_51_sram;
wire [0:3] mux_tree_tapbuf_size11_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_52_sram;
wire [0:3] mux_tree_tapbuf_size11_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_53_sram;
wire [0:3] mux_tree_tapbuf_size11_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_54_sram;
wire [0:3] mux_tree_tapbuf_size11_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_55_sram;
wire [0:3] mux_tree_tapbuf_size11_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_56_sram;
wire [0:3] mux_tree_tapbuf_size11_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_57_sram;
wire [0:3] mux_tree_tapbuf_size11_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_58_sram;
wire [0:3] mux_tree_tapbuf_size11_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_59_sram;
wire [0:3] mux_tree_tapbuf_size11_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_60_sram;
wire [0:3] mux_tree_tapbuf_size11_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_61_sram;
wire [0:3] mux_tree_tapbuf_size11_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_62_sram;
wire [0:3] mux_tree_tapbuf_size11_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_63_sram;
wire [0:3] mux_tree_tapbuf_size11_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_64_sram;
wire [0:3] mux_tree_tapbuf_size11_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_65_sram;
wire [0:3] mux_tree_tapbuf_size11_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_66_sram;
wire [0:3] mux_tree_tapbuf_size11_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_67_sram;
wire [0:3] mux_tree_tapbuf_size11_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_68_sram;
wire [0:3] mux_tree_tapbuf_size11_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_69_sram;
wire [0:3] mux_tree_tapbuf_size11_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_70_sram;
wire [0:3] mux_tree_tapbuf_size11_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_71_sram;
wire [0:3] mux_tree_tapbuf_size11_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_36_sram;
wire [0:3] mux_tree_tapbuf_size12_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_37_sram;
wire [0:3] mux_tree_tapbuf_size12_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_38_sram;
wire [0:3] mux_tree_tapbuf_size12_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_39_sram;
wire [0:3] mux_tree_tapbuf_size12_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_40_sram;
wire [0:3] mux_tree_tapbuf_size12_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_41_sram;
wire [0:3] mux_tree_tapbuf_size12_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_42_sram;
wire [0:3] mux_tree_tapbuf_size12_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_43_sram;
wire [0:3] mux_tree_tapbuf_size12_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_44_sram;
wire [0:3] mux_tree_tapbuf_size12_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_45_sram;
wire [0:3] mux_tree_tapbuf_size12_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_46_sram;
wire [0:3] mux_tree_tapbuf_size12_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_47_sram;
wire [0:3] mux_tree_tapbuf_size12_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_48_sram;
wire [0:3] mux_tree_tapbuf_size12_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_49_sram;
wire [0:3] mux_tree_tapbuf_size12_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_50_sram;
wire [0:3] mux_tree_tapbuf_size12_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_51_sram;
wire [0:3] mux_tree_tapbuf_size12_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_52_sram;
wire [0:3] mux_tree_tapbuf_size12_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_53_sram;
wire [0:3] mux_tree_tapbuf_size12_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_54_sram;
wire [0:3] mux_tree_tapbuf_size12_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_55_sram;
wire [0:3] mux_tree_tapbuf_size12_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_56_sram;
wire [0:3] mux_tree_tapbuf_size12_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_57_sram;
wire [0:3] mux_tree_tapbuf_size12_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_58_sram;
wire [0:3] mux_tree_tapbuf_size12_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_59_sram;
wire [0:3] mux_tree_tapbuf_size12_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_60_sram;
wire [0:3] mux_tree_tapbuf_size12_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_61_sram;
wire [0:3] mux_tree_tapbuf_size12_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_62_sram;
wire [0:3] mux_tree_tapbuf_size12_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_63_sram;
wire [0:3] mux_tree_tapbuf_size12_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_64_sram;
wire [0:3] mux_tree_tapbuf_size12_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_65_sram;
wire [0:3] mux_tree_tapbuf_size12_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_66_sram;
wire [0:3] mux_tree_tapbuf_size12_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_67_sram;
wire [0:3] mux_tree_tapbuf_size12_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_68_sram;
wire [0:3] mux_tree_tapbuf_size12_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_69_sram;
wire [0:3] mux_tree_tapbuf_size12_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_70_sram;
wire [0:3] mux_tree_tapbuf_size12_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_71_sram;
wire [0:3] mux_tree_tapbuf_size12_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_72_sram;
wire [0:3] mux_tree_tapbuf_size12_72_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_73_sram;
wire [0:3] mux_tree_tapbuf_size12_73_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_74_sram;
wire [0:3] mux_tree_tapbuf_size12_74_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_75_sram;
wire [0:3] mux_tree_tapbuf_size12_75_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_76_sram;
wire [0:3] mux_tree_tapbuf_size12_76_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_77_sram;
wire [0:3] mux_tree_tapbuf_size12_77_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_78_sram;
wire [0:3] mux_tree_tapbuf_size12_78_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_79_sram;
wire [0:3] mux_tree_tapbuf_size12_79_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_80_sram;
wire [0:3] mux_tree_tapbuf_size12_80_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_81_sram;
wire [0:3] mux_tree_tapbuf_size12_81_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_82_sram;
wire [0:3] mux_tree_tapbuf_size12_82_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_83_sram;
wire [0:3] mux_tree_tapbuf_size12_83_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_84_sram;
wire [0:3] mux_tree_tapbuf_size12_84_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_85_sram;
wire [0:3] mux_tree_tapbuf_size12_85_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_86_sram;
wire [0:3] mux_tree_tapbuf_size12_86_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_87_sram;
wire [0:3] mux_tree_tapbuf_size12_87_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_88_sram;
wire [0:3] mux_tree_tapbuf_size12_88_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_10_sram;
wire [0:3] mux_tree_tapbuf_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_11_sram;
wire [0:3] mux_tree_tapbuf_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_12_sram;
wire [0:3] mux_tree_tapbuf_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_13_sram;
wire [0:3] mux_tree_tapbuf_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_9_sram;
wire [0:3] mux_tree_tapbuf_size13_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size15_0_sram;
wire [0:3] mux_tree_tapbuf_size15_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_1_sram;
wire [0:3] mux_tree_tapbuf_size15_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_1_ccff_tail;
wire [0:4] mux_tree_tapbuf_size16_0_sram;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_10_sram;
wire [0:4] mux_tree_tapbuf_size16_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_11_sram;
wire [0:4] mux_tree_tapbuf_size16_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_12_sram;
wire [0:4] mux_tree_tapbuf_size16_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_13_sram;
wire [0:4] mux_tree_tapbuf_size16_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_14_sram;
wire [0:4] mux_tree_tapbuf_size16_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_15_sram;
wire [0:4] mux_tree_tapbuf_size16_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_16_sram;
wire [0:4] mux_tree_tapbuf_size16_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_17_sram;
wire [0:4] mux_tree_tapbuf_size16_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_18_sram;
wire [0:4] mux_tree_tapbuf_size16_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_19_sram;
wire [0:4] mux_tree_tapbuf_size16_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_1_sram;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_20_sram;
wire [0:4] mux_tree_tapbuf_size16_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_21_sram;
wire [0:4] mux_tree_tapbuf_size16_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_22_sram;
wire [0:4] mux_tree_tapbuf_size16_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_23_sram;
wire [0:4] mux_tree_tapbuf_size16_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_24_sram;
wire [0:4] mux_tree_tapbuf_size16_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_2_sram;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_3_sram;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_4_sram;
wire [0:4] mux_tree_tapbuf_size16_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_5_sram;
wire [0:4] mux_tree_tapbuf_size16_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_6_sram;
wire [0:4] mux_tree_tapbuf_size16_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_7_sram;
wire [0:4] mux_tree_tapbuf_size16_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_8_sram;
wire [0:4] mux_tree_tapbuf_size16_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_9_sram;
wire [0:4] mux_tree_tapbuf_size16_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size17_0_sram;
wire [0:4] mux_tree_tapbuf_size17_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_10_sram;
wire [0:4] mux_tree_tapbuf_size17_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_11_sram;
wire [0:4] mux_tree_tapbuf_size17_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_12_sram;
wire [0:4] mux_tree_tapbuf_size17_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_13_sram;
wire [0:4] mux_tree_tapbuf_size17_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_14_sram;
wire [0:4] mux_tree_tapbuf_size17_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_15_sram;
wire [0:4] mux_tree_tapbuf_size17_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_16_sram;
wire [0:4] mux_tree_tapbuf_size17_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_17_sram;
wire [0:4] mux_tree_tapbuf_size17_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_1_sram;
wire [0:4] mux_tree_tapbuf_size17_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_2_sram;
wire [0:4] mux_tree_tapbuf_size17_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_3_sram;
wire [0:4] mux_tree_tapbuf_size17_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_4_sram;
wire [0:4] mux_tree_tapbuf_size17_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_5_sram;
wire [0:4] mux_tree_tapbuf_size17_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_6_sram;
wire [0:4] mux_tree_tapbuf_size17_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_7_sram;
wire [0:4] mux_tree_tapbuf_size17_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_8_sram;
wire [0:4] mux_tree_tapbuf_size17_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_9_sram;
wire [0:4] mux_tree_tapbuf_size17_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size17_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size18_0_sram;
wire [0:4] mux_tree_tapbuf_size18_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_1_sram;
wire [0:4] mux_tree_tapbuf_size18_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_2_sram;
wire [0:4] mux_tree_tapbuf_size18_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size18_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_2_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_34_sram;
wire [0:2] mux_tree_tapbuf_size5_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_35_sram;
wire [0:2] mux_tree_tapbuf_size5_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_36_sram;
wire [0:2] mux_tree_tapbuf_size5_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_1_sram;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 571 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 572 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 575 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 576 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 579 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 580 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 583 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 584 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 587 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 588 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 591 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 592 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 595 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 596 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 599 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 600 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 603 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 604 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 607 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 608 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 611 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 612 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 615 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 616 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 619 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 620 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 623 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 624 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 627 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 628 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 631 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 632 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 635 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 636 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 639 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 640 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 643 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 644 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 647 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 648 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 651 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 652 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 655 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 656 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 659 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 663 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 667 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 671 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 675 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 679 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 683 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 687 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 691 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 695 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 699 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 703 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 707 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 711 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 713 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 715 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 717 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 719 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 721 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 723 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 725 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 727 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 729 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 731 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 733 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 735 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 737 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 739 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 741 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 743 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 745 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 747 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 749 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 751 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 753 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 755 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 757 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 759 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 761 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size17 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[1], chanx_right_in[50], chanx_right_in[99], chanx_right_in[148]}),
		.sram(mux_tree_tapbuf_size17_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_0_sram_inv[0:4]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size17 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[6], chanx_right_in[55], chanx_right_in[104], chanx_right_in[153]}),
		.sram(mux_tree_tapbuf_size17_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_1_sram_inv[0:4]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size17 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[7], chanx_right_in[56], chanx_right_in[105], chanx_right_in[154]}),
		.sram(mux_tree_tapbuf_size17_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_2_sram_inv[0:4]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size17 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[9], chanx_right_in[58], chanx_right_in[107], chanx_right_in[156]}),
		.sram(mux_tree_tapbuf_size17_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_3_sram_inv[0:4]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size17 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[12], chanx_right_in[61], chanx_right_in[110], chanx_right_in[159]}),
		.sram(mux_tree_tapbuf_size17_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_4_sram_inv[0:4]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size17 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[13], chanx_right_in[62], chanx_right_in[111], chanx_right_in[160]}),
		.sram(mux_tree_tapbuf_size17_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_5_sram_inv[0:4]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size17 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[15], chanx_right_in[64], chanx_right_in[113], chanx_right_in[162]}),
		.sram(mux_tree_tapbuf_size17_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_6_sram_inv[0:4]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size17 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[16], chanx_right_in[65], chanx_right_in[114], chanx_right_in[163]}),
		.sram(mux_tree_tapbuf_size17_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_7_sram_inv[0:4]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size17 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[17], chanx_right_in[66], chanx_right_in[115], chanx_right_in[164]}),
		.sram(mux_tree_tapbuf_size17_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_8_sram_inv[0:4]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size17 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[20], chanx_right_in[69], chanx_right_in[118], chanx_right_in[167]}),
		.sram(mux_tree_tapbuf_size17_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_9_sram_inv[0:4]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size17 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[22], chanx_right_in[71], chanx_right_in[120], chanx_right_in[169]}),
		.sram(mux_tree_tapbuf_size17_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_10_sram_inv[0:4]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size17 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[24], chanx_right_in[73], chanx_right_in[122], chanx_right_in[171]}),
		.sram(mux_tree_tapbuf_size17_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_11_sram_inv[0:4]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size17 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[28], chanx_right_in[77], chanx_right_in[126], chanx_right_in[175]}),
		.sram(mux_tree_tapbuf_size17_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_12_sram_inv[0:4]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size17 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[31], chanx_right_in[80], chanx_right_in[129], chanx_right_in[178]}),
		.sram(mux_tree_tapbuf_size17_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_13_sram_inv[0:4]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size17 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[34], chanx_right_in[83], chanx_right_in[132], chanx_right_in[181]}),
		.sram(mux_tree_tapbuf_size17_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_14_sram_inv[0:4]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size17 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[36], chanx_right_in[85], chanx_right_in[134], chanx_right_in[183]}),
		.sram(mux_tree_tapbuf_size17_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_15_sram_inv[0:4]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size17 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[42], chanx_right_in[91], chanx_right_in[140], chanx_right_in[189]}),
		.sram(mux_tree_tapbuf_size17_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_16_sram_inv[0:4]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size17 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[44], chanx_right_in[93], chanx_right_in[142], chanx_right_in[191]}),
		.sram(mux_tree_tapbuf_size17_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_17_sram_inv[0:4]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size17_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_0_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_1_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_2_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_3_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_4_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_5_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_6_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_7_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_8_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_9_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_10_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_11_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_12_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_13_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_14_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_15_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_16_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_17_sram_inv[0:4]));

	mux_tree_tapbuf_size16 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, chanx_right_in[2], chanx_right_in[51], chanx_right_in[100], chanx_right_in[149]}),
		.sram(mux_tree_tapbuf_size16_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_0_sram_inv[0:4]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size16 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[3], chanx_right_in[52], chanx_right_in[101], chanx_right_in[150]}),
		.sram(mux_tree_tapbuf_size16_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_1_sram_inv[0:4]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size16 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, chanx_right_in[5], chanx_right_in[54], chanx_right_in[103], chanx_right_in[152]}),
		.sram(mux_tree_tapbuf_size16_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_2_sram_inv[0:4]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size16 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[8], chanx_right_in[57], chanx_right_in[106], chanx_right_in[155]}),
		.sram(mux_tree_tapbuf_size16_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_3_sram_inv[0:4]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size16 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[10], chanx_right_in[59], chanx_right_in[108], chanx_right_in[157]}),
		.sram(mux_tree_tapbuf_size16_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_4_sram_inv[0:4]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size16 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, chanx_right_in[11], chanx_right_in[60], chanx_right_in[109], chanx_right_in[158]}),
		.sram(mux_tree_tapbuf_size16_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_5_sram_inv[0:4]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size16 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, chanx_right_in[14], chanx_right_in[63], chanx_right_in[112], chanx_right_in[161]}),
		.sram(mux_tree_tapbuf_size16_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_6_sram_inv[0:4]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size16 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[18], chanx_right_in[67], chanx_right_in[116], chanx_right_in[165]}),
		.sram(mux_tree_tapbuf_size16_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_7_sram_inv[0:4]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size16 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[19], chanx_right_in[68], chanx_right_in[117], chanx_right_in[166]}),
		.sram(mux_tree_tapbuf_size16_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_8_sram_inv[0:4]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size16 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[21], chanx_right_in[70], chanx_right_in[119], chanx_right_in[168]}),
		.sram(mux_tree_tapbuf_size16_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_9_sram_inv[0:4]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size16 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, chanx_right_in[23], chanx_right_in[72], chanx_right_in[121], chanx_right_in[170]}),
		.sram(mux_tree_tapbuf_size16_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_10_sram_inv[0:4]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size16 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[26], chanx_right_in[75], chanx_right_in[124], chanx_right_in[173]}),
		.sram(mux_tree_tapbuf_size16_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_11_sram_inv[0:4]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size16 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[27], chanx_right_in[76], chanx_right_in[125], chanx_right_in[174]}),
		.sram(mux_tree_tapbuf_size16_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_12_sram_inv[0:4]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size16 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, chanx_right_in[29], chanx_right_in[78], chanx_right_in[127], chanx_right_in[176]}),
		.sram(mux_tree_tapbuf_size16_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_13_sram_inv[0:4]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size16 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[30], chanx_right_in[79], chanx_right_in[128], chanx_right_in[177]}),
		.sram(mux_tree_tapbuf_size16_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_14_sram_inv[0:4]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size16 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, chanx_right_in[32], chanx_right_in[81], chanx_right_in[130], chanx_right_in[179]}),
		.sram(mux_tree_tapbuf_size16_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_15_sram_inv[0:4]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size16 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[35], chanx_right_in[84], chanx_right_in[133], chanx_right_in[182]}),
		.sram(mux_tree_tapbuf_size16_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_16_sram_inv[0:4]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size16 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[37], chanx_right_in[86], chanx_right_in[135], chanx_right_in[184]}),
		.sram(mux_tree_tapbuf_size16_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_17_sram_inv[0:4]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size16 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, chanx_right_in[38], chanx_right_in[87], chanx_right_in[136], chanx_right_in[185]}),
		.sram(mux_tree_tapbuf_size16_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_18_sram_inv[0:4]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size16 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[39], chanx_right_in[88], chanx_right_in[137], chanx_right_in[186]}),
		.sram(mux_tree_tapbuf_size16_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_19_sram_inv[0:4]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size16 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[40], chanx_right_in[89], chanx_right_in[138], chanx_right_in[187]}),
		.sram(mux_tree_tapbuf_size16_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_20_sram_inv[0:4]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size16 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[41], chanx_right_in[90], chanx_right_in[139], chanx_right_in[188]}),
		.sram(mux_tree_tapbuf_size16_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_21_sram_inv[0:4]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size16 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[43], chanx_right_in[92], chanx_right_in[141], chanx_right_in[190]}),
		.sram(mux_tree_tapbuf_size16_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_22_sram_inv[0:4]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size16 mux_top_track_352 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[45], chanx_right_in[94], chanx_right_in[143], chanx_right_in[192]}),
		.sram(mux_tree_tapbuf_size16_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_23_sram_inv[0:4]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size16 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[0], chanx_right_in[49], chanx_right_in[98], chanx_right_in[147]}),
		.sram(mux_tree_tapbuf_size16_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_24_sram_inv[0:4]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size16_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_0_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_1_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_2_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_3_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_4_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_5_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_6_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_7_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_8_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_9_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_10_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_11_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_12_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_13_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_14_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_15_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_16_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_17_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_18_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_19_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_20_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_21_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_22_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_23_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_24_sram_inv[0:4]));

	mux_tree_tapbuf_size18 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[4], chanx_right_in[53], chanx_right_in[102], chanx_right_in[151]}),
		.sram(mux_tree_tapbuf_size18_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_0_sram_inv[0:4]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size18 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[25], chanx_right_in[74], chanx_right_in[123], chanx_right_in[172]}),
		.sram(mux_tree_tapbuf_size18_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_1_sram_inv[0:4]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size18 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[33], chanx_right_in[82], chanx_right_in[131], chanx_right_in[180]}),
		.sram(mux_tree_tapbuf_size18_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_2_sram_inv[0:4]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size18_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_0_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_1_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_2_sram_inv[0:4]));

	mux_tree_tapbuf_size15 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[46], chanx_right_in[95], chanx_right_in[144]}),
		.sram(mux_tree_tapbuf_size15_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_0_sram_inv[0:3]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size15 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[47], chanx_right_in[96], chanx_right_in[145]}),
		.sram(mux_tree_tapbuf_size15_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_1_sram_inv[0:3]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size15_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_0_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_1_sram_inv[0:3]));

	mux_tree_tapbuf_size14 mux_top_track_376 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[48], chanx_right_in[97], chanx_right_in[146]}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size14_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size11 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size11 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size11 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size11 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size11 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size11 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size11 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size11 mux_right_track_52 (
		.in({chany_top_in[33], chany_top_in[103], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size11 mux_right_track_64 (
		.in({chany_top_in[41], chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size11 mux_right_track_70 (
		.in({chany_top_in[45], chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size11 mux_right_track_84 (
		.in({chany_top_in[54], chany_top_in[167], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_11_sram_inv[0:3]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size11 mux_right_track_88 (
		.in({chany_top_in[57], chany_top_in[175], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_12_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size11 mux_right_track_104 (
		.in({chany_top_in[68], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[185]}),
		.sram(mux_tree_tapbuf_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_13_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size11 mux_right_track_106 (
		.in({chany_top_in[69], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[184]}),
		.sram(mux_tree_tapbuf_size11_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_14_sram_inv[0:3]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size11 mux_right_track_142 (
		.in({chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[160]}),
		.sram(mux_tree_tapbuf_size11_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_15_sram_inv[0:3]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size11 mux_right_track_160 (
		.in({chany_top_in[105], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[148]}),
		.sram(mux_tree_tapbuf_size11_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_16_sram_inv[0:3]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size11 mux_right_track_164 (
		.in({chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[145]}),
		.sram(mux_tree_tapbuf_size11_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_17_sram_inv[0:3]),
		.out(chanx_right_out[82]));

	mux_tree_tapbuf_size11 mux_right_track_180 (
		.in({chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[134]}),
		.sram(mux_tree_tapbuf_size11_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_18_sram_inv[0:3]),
		.out(chanx_right_out[90]));

	mux_tree_tapbuf_size11 mux_right_track_182 (
		.in({chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[133]}),
		.sram(mux_tree_tapbuf_size11_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_19_sram_inv[0:3]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_size11 mux_right_track_184 (
		.in({chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[132]}),
		.sram(mux_tree_tapbuf_size11_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_20_sram_inv[0:3]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size11 mux_right_track_186 (
		.in({chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[130]}),
		.sram(mux_tree_tapbuf_size11_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_21_sram_inv[0:3]),
		.out(chanx_right_out[93]));

	mux_tree_tapbuf_size11 mux_right_track_196 (
		.in({chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[124]}),
		.sram(mux_tree_tapbuf_size11_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_22_sram_inv[0:3]),
		.out(chanx_right_out[98]));

	mux_tree_tapbuf_size11 mux_right_track_198 (
		.in({chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[122]}),
		.sram(mux_tree_tapbuf_size11_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_23_sram_inv[0:3]),
		.out(chanx_right_out[99]));

	mux_tree_tapbuf_size11 mux_right_track_200 (
		.in({chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[121]}),
		.sram(mux_tree_tapbuf_size11_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_24_sram_inv[0:3]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size11 mux_right_track_202 (
		.in({chany_top_in[133], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[120]}),
		.sram(mux_tree_tapbuf_size11_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_25_sram_inv[0:3]),
		.out(chanx_right_out[101]));

	mux_tree_tapbuf_size11 mux_right_track_204 (
		.in({chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[118]}),
		.sram(mux_tree_tapbuf_size11_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_26_sram_inv[0:3]),
		.out(chanx_right_out[102]));

	mux_tree_tapbuf_size11 mux_right_track_208 (
		.in({chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[116]}),
		.sram(mux_tree_tapbuf_size11_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_27_sram_inv[0:3]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size11 mux_right_track_214 (
		.in({chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[112]}),
		.sram(mux_tree_tapbuf_size11_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_28_sram_inv[0:3]),
		.out(chanx_right_out[107]));

	mux_tree_tapbuf_size11 mux_right_track_218 (
		.in({chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[109]}),
		.sram(mux_tree_tapbuf_size11_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_29_sram_inv[0:3]),
		.out(chanx_right_out[109]));

	mux_tree_tapbuf_size11 mux_right_track_220 (
		.in({chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[108]}),
		.sram(mux_tree_tapbuf_size11_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_30_sram_inv[0:3]),
		.out(chanx_right_out[110]));

	mux_tree_tapbuf_size11 mux_right_track_222 (
		.in({chany_top_in[146], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[106]}),
		.sram(mux_tree_tapbuf_size11_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_31_sram_inv[0:3]),
		.out(chanx_right_out[111]));

	mux_tree_tapbuf_size11 mux_right_track_226 (
		.in({chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[104]}),
		.sram(mux_tree_tapbuf_size11_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_32_sram_inv[0:3]),
		.out(chanx_right_out[113]));

	mux_tree_tapbuf_size11 mux_right_track_228 (
		.in({chany_top_in[150], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size11_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_33_sram_inv[0:3]),
		.out(chanx_right_out[114]));

	mux_tree_tapbuf_size11 mux_right_track_232 (
		.in({chany_top_in[153], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size11_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_34_sram_inv[0:3]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size11 mux_right_track_238 (
		.in({chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[96]}),
		.sram(mux_tree_tapbuf_size11_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_35_sram_inv[0:3]),
		.out(chanx_right_out[119]));

	mux_tree_tapbuf_size11 mux_right_track_240 (
		.in({chany_top_in[158], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[94]}),
		.sram(mux_tree_tapbuf_size11_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_36_sram_inv[0:3]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size11 mux_right_track_244 (
		.in({chany_top_in[161], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_size11_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_37_sram_inv[0:3]),
		.out(chanx_right_out[122]));

	mux_tree_tapbuf_size11 mux_right_track_246 (
		.in({chany_top_in[162], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size11_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_38_sram_inv[0:3]),
		.out(chanx_right_out[123]));

	mux_tree_tapbuf_size11 mux_right_track_248 (
		.in({chany_top_in[164], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_size11_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_39_sram_inv[0:3]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size11 mux_right_track_258 (
		.in({chany_top_in[170], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[82]}),
		.sram(mux_tree_tapbuf_size11_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_40_sram_inv[0:3]),
		.out(chanx_right_out[129]));

	mux_tree_tapbuf_size11 mux_right_track_262 (
		.in({chany_top_in[173], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[80]}),
		.sram(mux_tree_tapbuf_size11_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_41_sram_inv[0:3]),
		.out(chanx_right_out[131]));

	mux_tree_tapbuf_size11 mux_right_track_264 (
		.in({chany_top_in[174], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[78]}),
		.sram(mux_tree_tapbuf_size11_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_42_sram_inv[0:3]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size11 mux_right_track_266 (
		.in({chany_top_in[176], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size11_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_43_sram_inv[0:3]),
		.out(chanx_right_out[133]));

	mux_tree_tapbuf_size11 mux_right_track_280 (
		.in({chany_top_in[185], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_size11_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_44_sram_inv[0:3]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size11 mux_right_track_282 (
		.in({chany_top_in[186], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[66]}),
		.sram(mux_tree_tapbuf_size11_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_45_sram_inv[0:3]),
		.out(chanx_right_out[141]));

	mux_tree_tapbuf_size11 mux_right_track_284 (
		.in({chany_top_in[188], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_size11_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_46_sram_inv[0:3]),
		.out(chanx_right_out[142]));

	mux_tree_tapbuf_size11 mux_right_track_286 (
		.in({chany_top_in[189], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[64], chany_bottom_in[192]}),
		.sram(mux_tree_tapbuf_size11_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_47_sram_inv[0:3]),
		.out(chanx_right_out[143]));

	mux_tree_tapbuf_size11 mux_right_track_298 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[56], chany_bottom_in[171]}),
		.sram(mux_tree_tapbuf_size11_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_48_sram_inv[0:3]),
		.out(chanx_right_out[149]));

	mux_tree_tapbuf_size11 mux_right_track_300 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[54], chany_bottom_in[167]}),
		.sram(mux_tree_tapbuf_size11_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_49_sram_inv[0:3]),
		.out(chanx_right_out[150]));

	mux_tree_tapbuf_size11 mux_right_track_302 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[53], chany_bottom_in[163]}),
		.sram(mux_tree_tapbuf_size11_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_50_sram_inv[0:3]),
		.out(chanx_right_out[151]));

	mux_tree_tapbuf_size11 mux_right_track_306 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[50], chany_bottom_in[155]}),
		.sram(mux_tree_tapbuf_size11_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_51_sram_inv[0:3]),
		.out(chanx_right_out[153]));

	mux_tree_tapbuf_size11 mux_right_track_308 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[49], chany_bottom_in[151]}),
		.sram(mux_tree_tapbuf_size11_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_52_sram_inv[0:3]),
		.out(chanx_right_out[154]));

	mux_tree_tapbuf_size11 mux_right_track_318 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[42], chany_bottom_in[131]}),
		.sram(mux_tree_tapbuf_size11_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_53_sram_inv[0:3]),
		.out(chanx_right_out[159]));

	mux_tree_tapbuf_size11 mux_right_track_320 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[41], chany_bottom_in[127]}),
		.sram(mux_tree_tapbuf_size11_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_54_sram_inv[0:3]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size11 mux_right_track_324 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[38], chany_bottom_in[119]}),
		.sram(mux_tree_tapbuf_size11_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_55_sram_inv[0:3]),
		.out(chanx_right_out[162]));

	mux_tree_tapbuf_size11 mux_right_track_326 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[37], chany_bottom_in[115]}),
		.sram(mux_tree_tapbuf_size11_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_56_sram_inv[0:3]),
		.out(chanx_right_out[163]));

	mux_tree_tapbuf_size11 mux_right_track_328 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[36], chany_bottom_in[111]}),
		.sram(mux_tree_tapbuf_size11_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_57_sram_inv[0:3]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size11 mux_right_track_338 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[29], chany_bottom_in[91]}),
		.sram(mux_tree_tapbuf_size11_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_58_sram_inv[0:3]),
		.out(chanx_right_out[169]));

	mux_tree_tapbuf_size11 mux_right_track_342 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[26], chany_bottom_in[83]}),
		.sram(mux_tree_tapbuf_size11_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_59_sram_inv[0:3]),
		.out(chanx_right_out[171]));

	mux_tree_tapbuf_size11 mux_right_track_344 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[25], chany_bottom_in[79]}),
		.sram(mux_tree_tapbuf_size11_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_60_sram_inv[0:3]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size11 mux_right_track_346 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_size11_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_61_sram_inv[0:3]),
		.out(chanx_right_out[173]));

	mux_tree_tapbuf_size11 mux_right_track_348 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_size11_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_62_sram_inv[0:3]),
		.out(chanx_right_out[174]));

	mux_tree_tapbuf_size11 mux_right_track_350 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size11_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_63_sram_inv[0:3]),
		.out(chanx_right_out[175]));

	mux_tree_tapbuf_size11 mux_right_track_360 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size11_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_64_sram_inv[0:3]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size11 mux_right_track_362 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size11_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_65_sram_inv[0:3]),
		.out(chanx_right_out[181]));

	mux_tree_tapbuf_size11 mux_right_track_364 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size11_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_66_sram_inv[0:3]),
		.out(chanx_right_out[182]));

	mux_tree_tapbuf_size11 mux_right_track_366 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size11_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_67_sram_inv[0:3]),
		.out(chanx_right_out[183]));

	mux_tree_tapbuf_size11 mux_right_track_376 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size11_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_68_sram_inv[0:3]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size11 mux_right_track_378 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size11_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_69_sram_inv[0:3]),
		.out(chanx_right_out[189]));

	mux_tree_tapbuf_size11 mux_right_track_380 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size11_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_70_sram_inv[0:3]),
		.out(chanx_right_out[190]));

	mux_tree_tapbuf_size11 mux_right_track_382 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_size11_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_71_sram_inv[0:3]),
		.out(chanx_right_out[191]));

	mux_tree_tapbuf_size11_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_14_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_15_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_16_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_17_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_18_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_19_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_20_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_21_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_22_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_23_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_24_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_25_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_26_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_27_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_28_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_29_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_30_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_31_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_32_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_33_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_34_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_35_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_36_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_37_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_38_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_39_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_40_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_41_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_42_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_43_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_44_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_45_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_46_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_47_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_48_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_49_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_50_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_51_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_52_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_53_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_54_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_55_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_56_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_57_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_58_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_59_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_60_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_61_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_62_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_63_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_64_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_65_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_66_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_67_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_68_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_378 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_69_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_380 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_70_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_382 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_71_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size12 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size12 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size12 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size12 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size12 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size12 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size12 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size12 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size12 mux_right_track_40 (
		.in({chany_top_in[25], chany_top_in[79], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size12 mux_right_track_42 (
		.in({chany_top_in[26], chany_top_in[83], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size12 mux_right_track_46 (
		.in({chany_top_in[29], chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size12 mux_right_track_48 (
		.in({chany_top_in[30], chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size12 mux_right_track_50 (
		.in({chany_top_in[32], chany_top_in[99], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size12 mux_right_track_56 (
		.in({chany_top_in[36], chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size12 mux_right_track_58 (
		.in({chany_top_in[37], chany_top_in[115], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size12 mux_right_track_60 (
		.in({chany_top_in[38], chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size12 mux_right_track_62 (
		.in({chany_top_in[40], chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size12 mux_right_track_66 (
		.in({chany_top_in[42], chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size12 mux_right_track_68 (
		.in({chany_top_in[44], chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size12 mux_right_track_74 (
		.in({chany_top_in[48], chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size12 mux_right_track_76 (
		.in({chany_top_in[49], chany_top_in[151], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size12 mux_right_track_78 (
		.in({chany_top_in[50], chany_top_in[155], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size12 mux_right_track_80 (
		.in({chany_top_in[52], chany_top_in[159], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size12 mux_right_track_82 (
		.in({chany_top_in[53], chany_top_in[163], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size12 mux_right_track_86 (
		.in({chany_top_in[56], chany_top_in[171], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size12 mux_right_track_92 (
		.in({chany_top_in[60], chany_top_in[183], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size12 mux_right_track_94 (
		.in({chany_top_in[61], chany_top_in[187], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size12 mux_right_track_100 (
		.in({chany_top_in[65], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[188]}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size12 mux_right_track_102 (
		.in({chany_top_in[66], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[186]}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size12 mux_right_track_110 (
		.in({chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[181]}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size12 mux_right_track_112 (
		.in({chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[180]}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size12 mux_right_track_114 (
		.in({chany_top_in[74], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[178]}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size12 mux_right_track_116 (
		.in({chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[177]}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size12 mux_right_track_118 (
		.in({chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[176]}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size12 mux_right_track_120 (
		.in({chany_top_in[78], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[174]}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size12 mux_right_track_122 (
		.in({chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[173]}),
		.sram(mux_tree_tapbuf_size12_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_36_sram_inv[0:3]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size12 mux_right_track_128 (
		.in({chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[169]}),
		.sram(mux_tree_tapbuf_size12_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_37_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size12 mux_right_track_130 (
		.in({chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[168]}),
		.sram(mux_tree_tapbuf_size12_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_38_sram_inv[0:3]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size12 mux_right_track_132 (
		.in({chany_top_in[86], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[166]}),
		.sram(mux_tree_tapbuf_size12_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_39_sram_inv[0:3]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size12 mux_right_track_134 (
		.in({chany_top_in[88], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[165]}),
		.sram(mux_tree_tapbuf_size12_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_40_sram_inv[0:3]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size12 mux_right_track_136 (
		.in({chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[164]}),
		.sram(mux_tree_tapbuf_size12_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_41_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size12 mux_right_track_138 (
		.in({chany_top_in[90], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[162]}),
		.sram(mux_tree_tapbuf_size12_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_42_sram_inv[0:3]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size12 mux_right_track_140 (
		.in({chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[161]}),
		.sram(mux_tree_tapbuf_size12_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_43_sram_inv[0:3]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size12 mux_right_track_144 (
		.in({chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[158]}),
		.sram(mux_tree_tapbuf_size12_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_44_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size12 mux_right_track_146 (
		.in({chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[157]}),
		.sram(mux_tree_tapbuf_size12_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_45_sram_inv[0:3]),
		.out(chanx_right_out[73]));

	mux_tree_tapbuf_size12 mux_right_track_148 (
		.in({chany_top_in[97], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[156]}),
		.sram(mux_tree_tapbuf_size12_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_46_sram_inv[0:3]),
		.out(chanx_right_out[74]));

	mux_tree_tapbuf_size12 mux_right_track_150 (
		.in({chany_top_in[98], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[154]}),
		.sram(mux_tree_tapbuf_size12_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_47_sram_inv[0:3]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_size12 mux_right_track_152 (
		.in({chany_top_in[100], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[153]}),
		.sram(mux_tree_tapbuf_size12_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_48_sram_inv[0:3]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size12 mux_right_track_154 (
		.in({chany_top_in[101], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[152]}),
		.sram(mux_tree_tapbuf_size12_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_49_sram_inv[0:3]),
		.out(chanx_right_out[77]));

	mux_tree_tapbuf_size12 mux_right_track_156 (
		.in({chany_top_in[102], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[150]}),
		.sram(mux_tree_tapbuf_size12_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_50_sram_inv[0:3]),
		.out(chanx_right_out[78]));

	mux_tree_tapbuf_size12 mux_right_track_158 (
		.in({chany_top_in[104], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[149]}),
		.sram(mux_tree_tapbuf_size12_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_51_sram_inv[0:3]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_size12 mux_right_track_166 (
		.in({chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[144]}),
		.sram(mux_tree_tapbuf_size12_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_52_sram_inv[0:3]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_size12 mux_right_track_168 (
		.in({chany_top_in[110], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[142]}),
		.sram(mux_tree_tapbuf_size12_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_53_sram_inv[0:3]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size12 mux_right_track_170 (
		.in({chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[141]}),
		.sram(mux_tree_tapbuf_size12_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_54_sram_inv[0:3]),
		.out(chanx_right_out[85]));

	mux_tree_tapbuf_size12 mux_right_track_172 (
		.in({chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[140]}),
		.sram(mux_tree_tapbuf_size12_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_55_sram_inv[0:3]),
		.out(chanx_right_out[86]));

	mux_tree_tapbuf_size12 mux_right_track_174 (
		.in({chany_top_in[114], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[138]}),
		.sram(mux_tree_tapbuf_size12_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_56_sram_inv[0:3]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_size12 mux_right_track_176 (
		.in({chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[137]}),
		.sram(mux_tree_tapbuf_size12_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_57_sram_inv[0:3]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size12 mux_right_track_188 (
		.in({chany_top_in[124], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[129]}),
		.sram(mux_tree_tapbuf_size12_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_58_sram_inv[0:3]),
		.out(chanx_right_out[94]));

	mux_tree_tapbuf_size12 mux_right_track_192 (
		.in({chany_top_in[126], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[126]}),
		.sram(mux_tree_tapbuf_size12_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_59_sram_inv[0:3]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size12 mux_right_track_194 (
		.in({chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[125]}),
		.sram(mux_tree_tapbuf_size12_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_60_sram_inv[0:3]),
		.out(chanx_right_out[97]));

	mux_tree_tapbuf_size12 mux_right_track_206 (
		.in({chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[117]}),
		.sram(mux_tree_tapbuf_size12_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_61_sram_inv[0:3]),
		.out(chanx_right_out[103]));

	mux_tree_tapbuf_size12 mux_right_track_212 (
		.in({chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[113]}),
		.sram(mux_tree_tapbuf_size12_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_62_sram_inv[0:3]),
		.out(chanx_right_out[106]));

	mux_tree_tapbuf_size12 mux_right_track_216 (
		.in({chany_top_in[142], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[110]}),
		.sram(mux_tree_tapbuf_size12_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_63_sram_inv[0:3]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size12 mux_right_track_224 (
		.in({chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[105]}),
		.sram(mux_tree_tapbuf_size12_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_64_sram_inv[0:3]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size12 mux_right_track_234 (
		.in({chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size12_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_65_sram_inv[0:3]),
		.out(chanx_right_out[117]));

	mux_tree_tapbuf_size12 mux_right_track_236 (
		.in({chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[97]}),
		.sram(mux_tree_tapbuf_size12_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_66_sram_inv[0:3]),
		.out(chanx_right_out[118]));

	mux_tree_tapbuf_size12 mux_right_track_242 (
		.in({chany_top_in[160], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[93]}),
		.sram(mux_tree_tapbuf_size12_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_67_sram_inv[0:3]),
		.out(chanx_right_out[121]));

	mux_tree_tapbuf_size12 mux_right_track_252 (
		.in({chany_top_in[166], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_size12_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_68_sram_inv[0:3]),
		.out(chanx_right_out[126]));

	mux_tree_tapbuf_size12 mux_right_track_254 (
		.in({chany_top_in[168], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_size12_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_69_sram_inv[0:3]),
		.out(chanx_right_out[127]));

	mux_tree_tapbuf_size12 mux_right_track_256 (
		.in({chany_top_in[169], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[84]}),
		.sram(mux_tree_tapbuf_size12_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_70_sram_inv[0:3]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size12 mux_right_track_260 (
		.in({chany_top_in[172], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[81]}),
		.sram(mux_tree_tapbuf_size12_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_71_sram_inv[0:3]),
		.out(chanx_right_out[130]));

	mux_tree_tapbuf_size12 mux_right_track_272 (
		.in({chany_top_in[180], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_size12_72_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_72_sram_inv[0:3]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size12 mux_right_track_274 (
		.in({chany_top_in[181], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size12_73_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_73_sram_inv[0:3]),
		.out(chanx_right_out[137]));

	mux_tree_tapbuf_size12 mux_right_track_276 (
		.in({chany_top_in[182], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[70]}),
		.sram(mux_tree_tapbuf_size12_74_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_74_sram_inv[0:3]),
		.out(chanx_right_out[138]));

	mux_tree_tapbuf_size12 mux_right_track_278 (
		.in({chany_top_in[184], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_size12_75_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_75_sram_inv[0:3]),
		.out(chanx_right_out[139]));

	mux_tree_tapbuf_size12 mux_right_track_288 (
		.in({chany_top_in[190], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[62], chany_bottom_in[191]}),
		.sram(mux_tree_tapbuf_size12_76_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_76_sram_inv[0:3]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size12 mux_right_track_292 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[60], chany_bottom_in[183]}),
		.sram(mux_tree_tapbuf_size12_77_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_77_sram_inv[0:3]),
		.out(chanx_right_out[146]));

	mux_tree_tapbuf_size12 mux_right_track_294 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[58], chany_bottom_in[179]}),
		.sram(mux_tree_tapbuf_size12_78_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_78_sram_inv[0:3]),
		.out(chanx_right_out[147]));

	mux_tree_tapbuf_size12 mux_right_track_312 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[46], chany_bottom_in[143]}),
		.sram(mux_tree_tapbuf_size12_79_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_79_sram_inv[0:3]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size12 mux_right_track_316 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[44], chany_bottom_in[135]}),
		.sram(mux_tree_tapbuf_size12_80_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_80_sram_inv[0:3]),
		.out(chanx_right_out[158]));

	mux_tree_tapbuf_size12 mux_right_track_334 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[32], chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size12_81_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_81_sram_inv[0:3]),
		.out(chanx_right_out[167]));

	mux_tree_tapbuf_size12 mux_right_track_336 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[30], chany_bottom_in[95]}),
		.sram(mux_tree_tapbuf_size12_82_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_82_sram_inv[0:3]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size12 mux_right_track_352 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size12_83_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_83_sram_inv[0:3]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size12 mux_right_track_354 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size12_84_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_84_sram_inv[0:3]),
		.out(chanx_right_out[177]));

	mux_tree_tapbuf_size12 mux_right_track_356 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size12_85_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_85_sram_inv[0:3]),
		.out(chanx_right_out[178]));

	mux_tree_tapbuf_size12 mux_right_track_368 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size12_86_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_86_sram_inv[0:3]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size12 mux_right_track_372 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size12_87_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_87_sram_inv[0:3]),
		.out(chanx_right_out[186]));

	mux_tree_tapbuf_size12 mux_right_track_374 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size12_88_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_88_sram_inv[0:3]),
		.out(chanx_right_out[187]));

	mux_tree_tapbuf_size12_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_36_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_37_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_38_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_39_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_40_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_41_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_42_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_43_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_44_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_45_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_46_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_47_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_48_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_49_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_50_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_51_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_52_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_53_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_54_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_55_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_56_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_57_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_58_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_59_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_60_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_61_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_62_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_63_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_64_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_65_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_66_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_67_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_68_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_69_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_70_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_71_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_72_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_72_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_73_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_73_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_74_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_74_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_75_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_75_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_76_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_76_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_77_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_77_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_78_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_78_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_79_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_79_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_80_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_80_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_81_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_81_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_82_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_82_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_83_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_83_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_84_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_84_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_85_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_85_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_86_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_86_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_87_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_87_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_88_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_88_sram_inv[0:3]));

	mux_tree_tapbuf_size13 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size13 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size13 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size13 mux_right_track_54 (
		.in({chany_top_in[34], chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size13 mux_right_track_72 (
		.in({chany_top_in[46], chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size13 mux_right_track_90 (
		.in({chany_top_in[58], chany_top_in[179], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size13 mux_right_track_96 (
		.in({chany_top_in[62], chany_top_in[191], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[190]}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size13 mux_right_track_98 (
		.in({chany_top_in[64], chany_top_in[192], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[189]}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size13 mux_right_track_108 (
		.in({chany_top_in[70], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[182]}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size13 mux_right_track_126 (
		.in({chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[170]}),
		.sram(mux_tree_tapbuf_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_9_sram_inv[0:3]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size13 mux_right_track_162 (
		.in({chany_top_in[106], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[146]}),
		.sram(mux_tree_tapbuf_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_10_sram_inv[0:3]),
		.out(chanx_right_out[81]));

	mux_tree_tapbuf_size13 mux_right_track_296 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[57], chany_bottom_in[175]}),
		.sram(mux_tree_tapbuf_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_11_sram_inv[0:3]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size13 mux_right_track_314 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[45], chany_bottom_in[139]}),
		.sram(mux_tree_tapbuf_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_12_sram_inv[0:3]),
		.out(chanx_right_out[157]));

	mux_tree_tapbuf_size13 mux_right_track_332 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[33], chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_13_sram_inv[0:3]),
		.out(chanx_right_out[166]));

	mux_tree_tapbuf_size13_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_size10 mux_right_track_44 (
		.in({chany_top_in[28], chany_top_in[87], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size10 mux_right_track_124 (
		.in({chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[172]}),
		.sram(mux_tree_tapbuf_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_1_sram_inv[0:3]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size10 mux_right_track_178 (
		.in({chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[136]}),
		.sram(mux_tree_tapbuf_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_2_sram_inv[0:3]),
		.out(chanx_right_out[89]));

	mux_tree_tapbuf_size10 mux_right_track_190 (
		.in({chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[128]}),
		.sram(mux_tree_tapbuf_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_3_sram_inv[0:3]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_size10 mux_right_track_210 (
		.in({chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[114]}),
		.sram(mux_tree_tapbuf_size10_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_4_sram_inv[0:3]),
		.out(chanx_right_out[105]));

	mux_tree_tapbuf_size10 mux_right_track_230 (
		.in({chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size10_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_5_sram_inv[0:3]),
		.out(chanx_right_out[115]));

	mux_tree_tapbuf_size10 mux_right_track_268 (
		.in({chany_top_in[177], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[76]}),
		.sram(mux_tree_tapbuf_size10_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_6_sram_inv[0:3]),
		.out(chanx_right_out[134]));

	mux_tree_tapbuf_size10 mux_right_track_270 (
		.in({chany_top_in[178], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_size10_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_7_sram_inv[0:3]),
		.out(chanx_right_out[135]));

	mux_tree_tapbuf_size10 mux_right_track_290 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[61], chany_bottom_in[187]}),
		.sram(mux_tree_tapbuf_size10_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_8_sram_inv[0:3]),
		.out(chanx_right_out[145]));

	mux_tree_tapbuf_size10 mux_right_track_304 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[52], chany_bottom_in[159]}),
		.sram(mux_tree_tapbuf_size10_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_9_sram_inv[0:3]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size10 mux_right_track_310 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[48], chany_bottom_in[147]}),
		.sram(mux_tree_tapbuf_size10_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_10_sram_inv[0:3]),
		.out(chanx_right_out[155]));

	mux_tree_tapbuf_size10 mux_right_track_322 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[40], chany_bottom_in[123]}),
		.sram(mux_tree_tapbuf_size10_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_11_sram_inv[0:3]),
		.out(chanx_right_out[161]));

	mux_tree_tapbuf_size10 mux_right_track_330 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[34], chany_bottom_in[107]}),
		.sram(mux_tree_tapbuf_size10_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_12_sram_inv[0:3]),
		.out(chanx_right_out[165]));

	mux_tree_tapbuf_size10 mux_right_track_340 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[28], chany_bottom_in[87]}),
		.sram(mux_tree_tapbuf_size10_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_13_sram_inv[0:3]),
		.out(chanx_right_out[170]));

	mux_tree_tapbuf_size10 mux_right_track_358 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size10_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_14_sram_inv[0:3]),
		.out(chanx_right_out[179]));

	mux_tree_tapbuf_size10 mux_right_track_370 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size10_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_15_sram_inv[0:3]),
		.out(chanx_right_out[185]));

	mux_tree_tapbuf_size10_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_4_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_5_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_6_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_7_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_8_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_9_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_10_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_11_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_12_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_13_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_14_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_15_sram_inv[0:3]));

	mux_tree_tapbuf_size9 mux_right_track_250 (
		.in({chany_top_in[165], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chanx_right_out[125]));

	mux_tree_tapbuf_size9 mux_right_track_384 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_1_sram_inv[0:3]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size9_mem mem_right_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_size5 mux_bottom_track_1 (
		.in({chanx_right_in[47], chanx_right_in[96], chanx_right_in[145], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size5 mux_bottom_track_9 (
		.in({chanx_right_in[46], chanx_right_in[95], chanx_right_in[144], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size5 mux_bottom_track_65 (
		.in({chanx_right_in[39], chanx_right_in[88], chanx_right_in[137], chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size5 mux_bottom_track_81 (
		.in({chanx_right_in[37], chanx_right_in[86], chanx_right_in[135], chanx_right_in[184], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size5 mux_bottom_track_89 (
		.in({chanx_right_in[36], chanx_right_in[85], chanx_right_in[134], chanx_right_in[183], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size5 mux_bottom_track_97 (
		.in({chanx_right_in[35], chanx_right_in[84], chanx_right_in[133], chanx_right_in[182], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size5 mux_bottom_track_105 (
		.in({chanx_right_in[34], chanx_right_in[83], chanx_right_in[132], chanx_right_in[181], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size5 mux_bottom_track_113 (
		.in({chanx_right_in[33], chanx_right_in[82], chanx_right_in[131], chanx_right_in[180], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size5 mux_bottom_track_121 (
		.in({chanx_right_in[32], chanx_right_in[81], chanx_right_in[130], chanx_right_in[179], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size5 mux_bottom_track_129 (
		.in({chanx_right_in[31], chanx_right_in[80], chanx_right_in[129], chanx_right_in[178], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size5 mux_bottom_track_137 (
		.in({chanx_right_in[30], chanx_right_in[79], chanx_right_in[128], chanx_right_in[177], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size5 mux_bottom_track_153 (
		.in({chanx_right_in[28], chanx_right_in[77], chanx_right_in[126], chanx_right_in[175], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size5 mux_bottom_track_161 (
		.in({chanx_right_in[27], chanx_right_in[76], chanx_right_in[125], chanx_right_in[174], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size5 mux_bottom_track_169 (
		.in({chanx_right_in[26], chanx_right_in[75], chanx_right_in[124], chanx_right_in[173], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size5 mux_bottom_track_177 (
		.in({chanx_right_in[25], chanx_right_in[74], chanx_right_in[123], chanx_right_in[172], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size5 mux_bottom_track_185 (
		.in({chanx_right_in[24], chanx_right_in[73], chanx_right_in[122], chanx_right_in[171], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size5 mux_bottom_track_193 (
		.in({chanx_right_in[23], chanx_right_in[72], chanx_right_in[121], chanx_right_in[170], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size5 mux_bottom_track_201 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[120], chanx_right_in[169], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size5 mux_bottom_track_209 (
		.in({chanx_right_in[21], chanx_right_in[70], chanx_right_in[119], chanx_right_in[168], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size5 mux_bottom_track_225 (
		.in({chanx_right_in[19], chanx_right_in[68], chanx_right_in[117], chanx_right_in[166], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size5 mux_bottom_track_233 (
		.in({chanx_right_in[18], chanx_right_in[67], chanx_right_in[116], chanx_right_in[165], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size5 mux_bottom_track_241 (
		.in({chanx_right_in[17], chanx_right_in[66], chanx_right_in[115], chanx_right_in[164], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size5 mux_bottom_track_249 (
		.in({chanx_right_in[16], chanx_right_in[65], chanx_right_in[114], chanx_right_in[163], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size5 mux_bottom_track_257 (
		.in({chanx_right_in[15], chanx_right_in[64], chanx_right_in[113], chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size5 mux_bottom_track_265 (
		.in({chanx_right_in[14], chanx_right_in[63], chanx_right_in[112], chanx_right_in[161], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size5 mux_bottom_track_273 (
		.in({chanx_right_in[13], chanx_right_in[62], chanx_right_in[111], chanx_right_in[160], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size5 mux_bottom_track_281 (
		.in({chanx_right_in[12], chanx_right_in[61], chanx_right_in[110], chanx_right_in[159], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size5 mux_bottom_track_297 (
		.in({chanx_right_in[10], chanx_right_in[59], chanx_right_in[108], chanx_right_in[157], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size5 mux_bottom_track_305 (
		.in({chanx_right_in[9], chanx_right_in[58], chanx_right_in[107], chanx_right_in[156], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size5 mux_bottom_track_313 (
		.in({chanx_right_in[8], chanx_right_in[57], chanx_right_in[106], chanx_right_in[155], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size5 mux_bottom_track_321 (
		.in({chanx_right_in[7], chanx_right_in[56], chanx_right_in[105], chanx_right_in[154], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size5 mux_bottom_track_329 (
		.in({chanx_right_in[6], chanx_right_in[55], chanx_right_in[104], chanx_right_in[153], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size5 mux_bottom_track_337 (
		.in({chanx_right_in[5], chanx_right_in[54], chanx_right_in[103], chanx_right_in[152], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size5 mux_bottom_track_345 (
		.in({chanx_right_in[4], chanx_right_in[53], chanx_right_in[102], chanx_right_in[151], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size5 mux_bottom_track_353 (
		.in({chanx_right_in[3], chanx_right_in[52], chanx_right_in[101], chanx_right_in[150], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_34_sram_inv[0:2]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size5 mux_bottom_track_369 (
		.in({chanx_right_in[1], chanx_right_in[50], chanx_right_in[99], chanx_right_in[148], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_35_sram_inv[0:2]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size5 mux_bottom_track_377 (
		.in({chanx_right_in[0], chanx_right_in[49], chanx_right_in[98], chanx_right_in[147], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_36_sram_inv[0:2]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_34_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_35_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_36_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_bottom_track_17 (
		.in({chanx_right_in[45], chanx_right_in[94], chanx_right_in[143], chanx_right_in[192], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size6 mux_bottom_track_25 (
		.in({chanx_right_in[44], chanx_right_in[93], chanx_right_in[142], chanx_right_in[191], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size6 mux_bottom_track_33 (
		.in({chanx_right_in[43], chanx_right_in[92], chanx_right_in[141], chanx_right_in[190], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size6 mux_bottom_track_41 (
		.in({chanx_right_in[42], chanx_right_in[91], chanx_right_in[140], chanx_right_in[189], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size6 mux_bottom_track_49 (
		.in({chanx_right_in[41], chanx_right_in[90], chanx_right_in[139], chanx_right_in[188], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_57 (
		.in({chanx_right_in[40], chanx_right_in[89], chanx_right_in[138], chanx_right_in[187], bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size6 mux_bottom_track_73 (
		.in({chanx_right_in[38], chanx_right_in[87], chanx_right_in[136], chanx_right_in[185], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size6 mux_bottom_track_145 (
		.in({chanx_right_in[29], chanx_right_in[78], chanx_right_in[127], chanx_right_in[176], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size6 mux_bottom_track_217 (
		.in({chanx_right_in[20], chanx_right_in[69], chanx_right_in[118], chanx_right_in[167], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size6 mux_bottom_track_289 (
		.in({chanx_right_in[11], chanx_right_in[60], chanx_right_in[109], chanx_right_in[158], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size6 mux_bottom_track_361 (
		.in({chanx_right_in[2], chanx_right_in[51], chanx_right_in[100], chanx_right_in[149], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_bottom_track_385 (
		.in({chanx_right_in[48], chanx_right_in[97], chanx_right_in[146], bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_bottom_out[192]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_0__1_ -----

//----- Default net type -----
`default_nettype wire



