//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for physical tile: router]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul 21 19:29:39 2024
//-------------------------------------------
// ----- BEGIN Grid Verilog module: grid_router -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for grid_router -----
module grid_router(clk,
                   set,
                   reset,
                   prog_clk,
                   top_width_0_height_0_subtile_0__pin_rst__0_,
                   top_width_0_height_0_subtile_0__pin_my_ypos_1_,
                   top_width_0_height_0_subtile_0__pin_idata_0_3_,
                   top_width_0_height_0_subtile_0__pin_idata_0_7_,
                   top_width_0_height_0_subtile_0__pin_idata_0_11_,
                   top_width_0_height_0_subtile_0__pin_idata_0_15_,
                   top_width_0_height_0_subtile_0__pin_idata_0_19_,
                   top_width_0_height_0_subtile_0__pin_idata_0_23_,
                   top_width_0_height_0_subtile_0__pin_idata_0_27_,
                   top_width_0_height_0_subtile_0__pin_idata_0_31_,
                   top_width_0_height_0_subtile_0__pin_idata_1_0_,
                   top_width_0_height_0_subtile_0__pin_idata_1_4_,
                   top_width_0_height_0_subtile_0__pin_idata_1_8_,
                   top_width_0_height_0_subtile_0__pin_idata_1_12_,
                   top_width_0_height_0_subtile_0__pin_idata_1_16_,
                   top_width_0_height_0_subtile_0__pin_idata_1_20_,
                   top_width_0_height_0_subtile_0__pin_idata_1_24_,
                   top_width_0_height_0_subtile_0__pin_idata_1_28_,
                   top_width_0_height_0_subtile_0__pin_idata_1_32_,
                   top_width_0_height_0_subtile_0__pin_idata_2_1_,
                   top_width_0_height_0_subtile_0__pin_idata_2_5_,
                   top_width_0_height_0_subtile_0__pin_idata_2_9_,
                   top_width_0_height_0_subtile_0__pin_idata_2_13_,
                   top_width_0_height_0_subtile_0__pin_idata_2_17_,
                   top_width_0_height_0_subtile_0__pin_idata_2_21_,
                   top_width_0_height_0_subtile_0__pin_idata_2_25_,
                   top_width_0_height_0_subtile_0__pin_idata_2_29_,
                   top_width_0_height_0_subtile_0__pin_idata_2_33_,
                   top_width_0_height_0_subtile_0__pin_idata_3_2_,
                   top_width_0_height_0_subtile_0__pin_idata_3_6_,
                   top_width_0_height_0_subtile_0__pin_idata_3_10_,
                   top_width_0_height_0_subtile_0__pin_idata_3_14_,
                   top_width_0_height_0_subtile_0__pin_idata_3_18_,
                   top_width_0_height_0_subtile_0__pin_idata_3_22_,
                   top_width_0_height_0_subtile_0__pin_idata_3_26_,
                   top_width_0_height_0_subtile_0__pin_idata_3_30_,
                   top_width_0_height_0_subtile_0__pin_idata_3_34_,
                   top_width_0_height_0_subtile_0__pin_idata_4_3_,
                   top_width_0_height_0_subtile_0__pin_idata_4_7_,
                   top_width_0_height_0_subtile_0__pin_idata_4_11_,
                   top_width_0_height_0_subtile_0__pin_idata_4_15_,
                   top_width_0_height_0_subtile_0__pin_idata_4_19_,
                   top_width_0_height_0_subtile_0__pin_idata_4_23_,
                   top_width_0_height_0_subtile_0__pin_idata_4_27_,
                   top_width_0_height_0_subtile_0__pin_idata_4_31_,
                   top_width_0_height_0_subtile_0__pin_ivalid_0_0_,
                   top_width_0_height_0_subtile_0__pin_ivalid_4_0_,
                   top_width_0_height_0_subtile_0__pin_ivch_3_0_,
                   top_width_0_height_0_subtile_0__pin_iack_1_0_,
                   top_width_0_height_0_subtile_0__pin_iack_3_0_,
                   top_width_0_height_0_subtile_0__pin_ilck_0_0_,
                   top_width_0_height_0_subtile_0__pin_ilck_2_0_,
                   top_width_0_height_0_subtile_0__pin_ilck_4_0_,
                   right_width_0_height_0_subtile_0__pin_my_xpos_0_,
                   right_width_0_height_0_subtile_0__pin_idata_0_0_,
                   right_width_0_height_0_subtile_0__pin_idata_0_4_,
                   right_width_0_height_0_subtile_0__pin_idata_0_8_,
                   right_width_0_height_0_subtile_0__pin_idata_0_12_,
                   right_width_0_height_0_subtile_0__pin_idata_0_16_,
                   right_width_0_height_0_subtile_0__pin_idata_0_20_,
                   right_width_0_height_0_subtile_0__pin_idata_0_24_,
                   right_width_0_height_0_subtile_0__pin_idata_0_28_,
                   right_width_0_height_0_subtile_0__pin_idata_0_32_,
                   right_width_0_height_0_subtile_0__pin_idata_1_1_,
                   right_width_0_height_0_subtile_0__pin_idata_1_5_,
                   right_width_0_height_0_subtile_0__pin_idata_1_9_,
                   right_width_0_height_0_subtile_0__pin_idata_1_13_,
                   right_width_0_height_0_subtile_0__pin_idata_1_17_,
                   right_width_0_height_0_subtile_0__pin_idata_1_21_,
                   right_width_0_height_0_subtile_0__pin_idata_1_25_,
                   right_width_0_height_0_subtile_0__pin_idata_1_29_,
                   right_width_0_height_0_subtile_0__pin_idata_1_33_,
                   right_width_0_height_0_subtile_0__pin_idata_2_2_,
                   right_width_0_height_0_subtile_0__pin_idata_2_6_,
                   right_width_0_height_0_subtile_0__pin_idata_2_10_,
                   right_width_0_height_0_subtile_0__pin_idata_2_14_,
                   right_width_0_height_0_subtile_0__pin_idata_2_18_,
                   right_width_0_height_0_subtile_0__pin_idata_2_22_,
                   right_width_0_height_0_subtile_0__pin_idata_2_26_,
                   right_width_0_height_0_subtile_0__pin_idata_2_30_,
                   right_width_0_height_0_subtile_0__pin_idata_2_34_,
                   right_width_0_height_0_subtile_0__pin_idata_3_3_,
                   right_width_0_height_0_subtile_0__pin_idata_3_7_,
                   right_width_0_height_0_subtile_0__pin_idata_3_11_,
                   right_width_0_height_0_subtile_0__pin_idata_3_15_,
                   right_width_0_height_0_subtile_0__pin_idata_3_19_,
                   right_width_0_height_0_subtile_0__pin_idata_3_23_,
                   right_width_0_height_0_subtile_0__pin_idata_3_27_,
                   right_width_0_height_0_subtile_0__pin_idata_3_31_,
                   right_width_0_height_0_subtile_0__pin_idata_4_0_,
                   right_width_0_height_0_subtile_0__pin_idata_4_4_,
                   right_width_0_height_0_subtile_0__pin_idata_4_8_,
                   right_width_0_height_0_subtile_0__pin_idata_4_12_,
                   right_width_0_height_0_subtile_0__pin_idata_4_16_,
                   right_width_0_height_0_subtile_0__pin_idata_4_20_,
                   right_width_0_height_0_subtile_0__pin_idata_4_24_,
                   right_width_0_height_0_subtile_0__pin_idata_4_28_,
                   right_width_0_height_0_subtile_0__pin_idata_4_32_,
                   right_width_0_height_0_subtile_0__pin_ivalid_1_0_,
                   right_width_0_height_0_subtile_0__pin_ivch_0_0_,
                   right_width_0_height_0_subtile_0__pin_ivch_4_0_,
                   right_width_0_height_0_subtile_0__pin_iack_1_1_,
                   right_width_0_height_0_subtile_0__pin_iack_3_1_,
                   right_width_0_height_0_subtile_0__pin_ilck_0_1_,
                   right_width_0_height_0_subtile_0__pin_ilck_2_1_,
                   right_width_0_height_0_subtile_0__pin_ilck_4_1_,
                   right_width_0_height_0_subtile_0__pin_clk_0_,
                   bottom_width_0_height_0_subtile_0__pin_my_xpos_1_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_1_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_5_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_9_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_13_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_17_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_21_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_25_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_29_,
                   bottom_width_0_height_0_subtile_0__pin_idata_0_33_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_2_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_6_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_10_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_14_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_18_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_22_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_26_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_30_,
                   bottom_width_0_height_0_subtile_0__pin_idata_1_34_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_3_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_7_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_11_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_15_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_19_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_23_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_27_,
                   bottom_width_0_height_0_subtile_0__pin_idata_2_31_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_0_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_4_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_8_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_12_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_16_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_20_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_24_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_28_,
                   bottom_width_0_height_0_subtile_0__pin_idata_3_32_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_1_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_5_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_9_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_13_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_17_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_21_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_25_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_29_,
                   bottom_width_0_height_0_subtile_0__pin_idata_4_33_,
                   bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_,
                   bottom_width_0_height_0_subtile_0__pin_ivch_1_0_,
                   bottom_width_0_height_0_subtile_0__pin_iack_0_0_,
                   bottom_width_0_height_0_subtile_0__pin_iack_2_0_,
                   bottom_width_0_height_0_subtile_0__pin_iack_4_0_,
                   bottom_width_0_height_0_subtile_0__pin_ilck_1_0_,
                   bottom_width_0_height_0_subtile_0__pin_ilck_3_0_,
                   left_width_0_height_0_subtile_0__pin_my_ypos_0_,
                   left_width_0_height_0_subtile_0__pin_idata_0_2_,
                   left_width_0_height_0_subtile_0__pin_idata_0_6_,
                   left_width_0_height_0_subtile_0__pin_idata_0_10_,
                   left_width_0_height_0_subtile_0__pin_idata_0_14_,
                   left_width_0_height_0_subtile_0__pin_idata_0_18_,
                   left_width_0_height_0_subtile_0__pin_idata_0_22_,
                   left_width_0_height_0_subtile_0__pin_idata_0_26_,
                   left_width_0_height_0_subtile_0__pin_idata_0_30_,
                   left_width_0_height_0_subtile_0__pin_idata_0_34_,
                   left_width_0_height_0_subtile_0__pin_idata_1_3_,
                   left_width_0_height_0_subtile_0__pin_idata_1_7_,
                   left_width_0_height_0_subtile_0__pin_idata_1_11_,
                   left_width_0_height_0_subtile_0__pin_idata_1_15_,
                   left_width_0_height_0_subtile_0__pin_idata_1_19_,
                   left_width_0_height_0_subtile_0__pin_idata_1_23_,
                   left_width_0_height_0_subtile_0__pin_idata_1_27_,
                   left_width_0_height_0_subtile_0__pin_idata_1_31_,
                   left_width_0_height_0_subtile_0__pin_idata_2_0_,
                   left_width_0_height_0_subtile_0__pin_idata_2_4_,
                   left_width_0_height_0_subtile_0__pin_idata_2_8_,
                   left_width_0_height_0_subtile_0__pin_idata_2_12_,
                   left_width_0_height_0_subtile_0__pin_idata_2_16_,
                   left_width_0_height_0_subtile_0__pin_idata_2_20_,
                   left_width_0_height_0_subtile_0__pin_idata_2_24_,
                   left_width_0_height_0_subtile_0__pin_idata_2_28_,
                   left_width_0_height_0_subtile_0__pin_idata_2_32_,
                   left_width_0_height_0_subtile_0__pin_idata_3_1_,
                   left_width_0_height_0_subtile_0__pin_idata_3_5_,
                   left_width_0_height_0_subtile_0__pin_idata_3_9_,
                   left_width_0_height_0_subtile_0__pin_idata_3_13_,
                   left_width_0_height_0_subtile_0__pin_idata_3_17_,
                   left_width_0_height_0_subtile_0__pin_idata_3_21_,
                   left_width_0_height_0_subtile_0__pin_idata_3_25_,
                   left_width_0_height_0_subtile_0__pin_idata_3_29_,
                   left_width_0_height_0_subtile_0__pin_idata_3_33_,
                   left_width_0_height_0_subtile_0__pin_idata_4_2_,
                   left_width_0_height_0_subtile_0__pin_idata_4_6_,
                   left_width_0_height_0_subtile_0__pin_idata_4_10_,
                   left_width_0_height_0_subtile_0__pin_idata_4_14_,
                   left_width_0_height_0_subtile_0__pin_idata_4_18_,
                   left_width_0_height_0_subtile_0__pin_idata_4_22_,
                   left_width_0_height_0_subtile_0__pin_idata_4_26_,
                   left_width_0_height_0_subtile_0__pin_idata_4_30_,
                   left_width_0_height_0_subtile_0__pin_idata_4_34_,
                   left_width_0_height_0_subtile_0__pin_ivalid_3_0_,
                   left_width_0_height_0_subtile_0__pin_ivch_2_0_,
                   left_width_0_height_0_subtile_0__pin_iack_0_1_,
                   left_width_0_height_0_subtile_0__pin_iack_2_1_,
                   left_width_0_height_0_subtile_0__pin_iack_4_1_,
                   left_width_0_height_0_subtile_0__pin_ilck_1_1_,
                   left_width_0_height_0_subtile_0__pin_ilck_3_1_,
                   ccff_head,
                   top_width_0_height_0_subtile_0__pin_odata_0_2_,
                   top_width_0_height_0_subtile_0__pin_odata_0_6_,
                   top_width_0_height_0_subtile_0__pin_odata_0_10_,
                   top_width_0_height_0_subtile_0__pin_odata_0_14_,
                   top_width_0_height_0_subtile_0__pin_odata_0_18_,
                   top_width_0_height_0_subtile_0__pin_odata_0_22_,
                   top_width_0_height_0_subtile_0__pin_odata_0_26_,
                   top_width_0_height_0_subtile_0__pin_odata_0_30_,
                   top_width_0_height_0_subtile_0__pin_odata_0_34_,
                   top_width_0_height_0_subtile_0__pin_odata_1_3_,
                   top_width_0_height_0_subtile_0__pin_odata_1_7_,
                   top_width_0_height_0_subtile_0__pin_odata_1_11_,
                   top_width_0_height_0_subtile_0__pin_odata_1_15_,
                   top_width_0_height_0_subtile_0__pin_odata_1_19_,
                   top_width_0_height_0_subtile_0__pin_odata_1_23_,
                   top_width_0_height_0_subtile_0__pin_odata_1_27_,
                   top_width_0_height_0_subtile_0__pin_odata_1_31_,
                   top_width_0_height_0_subtile_0__pin_odata_2_0_,
                   top_width_0_height_0_subtile_0__pin_odata_2_4_,
                   top_width_0_height_0_subtile_0__pin_odata_2_8_,
                   top_width_0_height_0_subtile_0__pin_odata_2_12_,
                   top_width_0_height_0_subtile_0__pin_odata_2_16_,
                   top_width_0_height_0_subtile_0__pin_odata_2_20_,
                   top_width_0_height_0_subtile_0__pin_odata_2_24_,
                   top_width_0_height_0_subtile_0__pin_odata_2_28_,
                   top_width_0_height_0_subtile_0__pin_odata_2_32_,
                   top_width_0_height_0_subtile_0__pin_odata_3_1_,
                   top_width_0_height_0_subtile_0__pin_odata_3_5_,
                   top_width_0_height_0_subtile_0__pin_odata_3_9_,
                   top_width_0_height_0_subtile_0__pin_odata_3_13_,
                   top_width_0_height_0_subtile_0__pin_odata_3_17_,
                   top_width_0_height_0_subtile_0__pin_odata_3_21_,
                   top_width_0_height_0_subtile_0__pin_odata_3_25_,
                   top_width_0_height_0_subtile_0__pin_odata_3_29_,
                   top_width_0_height_0_subtile_0__pin_odata_3_33_,
                   top_width_0_height_0_subtile_0__pin_odata_4_2_,
                   top_width_0_height_0_subtile_0__pin_odata_4_6_,
                   top_width_0_height_0_subtile_0__pin_odata_4_10_,
                   top_width_0_height_0_subtile_0__pin_odata_4_14_,
                   top_width_0_height_0_subtile_0__pin_odata_4_18_,
                   top_width_0_height_0_subtile_0__pin_odata_4_22_,
                   top_width_0_height_0_subtile_0__pin_odata_4_26_,
                   top_width_0_height_0_subtile_0__pin_odata_4_30_,
                   top_width_0_height_0_subtile_0__pin_odata_4_34_,
                   top_width_0_height_0_subtile_0__pin_ovalid_3_0_,
                   top_width_0_height_0_subtile_0__pin_ovch_2_0_,
                   top_width_0_height_0_subtile_0__pin_oack_0_1_,
                   top_width_0_height_0_subtile_0__pin_oack_2_1_,
                   top_width_0_height_0_subtile_0__pin_oack_4_1_,
                   top_width_0_height_0_subtile_0__pin_ordy_1_1_,
                   top_width_0_height_0_subtile_0__pin_ordy_3_1_,
                   top_width_0_height_0_subtile_0__pin_olck_0_1_,
                   top_width_0_height_0_subtile_0__pin_olck_2_1_,
                   top_width_0_height_0_subtile_0__pin_olck_4_1_,
                   right_width_0_height_0_subtile_0__pin_odata_0_3_,
                   right_width_0_height_0_subtile_0__pin_odata_0_7_,
                   right_width_0_height_0_subtile_0__pin_odata_0_11_,
                   right_width_0_height_0_subtile_0__pin_odata_0_15_,
                   right_width_0_height_0_subtile_0__pin_odata_0_19_,
                   right_width_0_height_0_subtile_0__pin_odata_0_23_,
                   right_width_0_height_0_subtile_0__pin_odata_0_27_,
                   right_width_0_height_0_subtile_0__pin_odata_0_31_,
                   right_width_0_height_0_subtile_0__pin_odata_1_0_,
                   right_width_0_height_0_subtile_0__pin_odata_1_4_,
                   right_width_0_height_0_subtile_0__pin_odata_1_8_,
                   right_width_0_height_0_subtile_0__pin_odata_1_12_,
                   right_width_0_height_0_subtile_0__pin_odata_1_16_,
                   right_width_0_height_0_subtile_0__pin_odata_1_20_,
                   right_width_0_height_0_subtile_0__pin_odata_1_24_,
                   right_width_0_height_0_subtile_0__pin_odata_1_28_,
                   right_width_0_height_0_subtile_0__pin_odata_1_32_,
                   right_width_0_height_0_subtile_0__pin_odata_2_1_,
                   right_width_0_height_0_subtile_0__pin_odata_2_5_,
                   right_width_0_height_0_subtile_0__pin_odata_2_9_,
                   right_width_0_height_0_subtile_0__pin_odata_2_13_,
                   right_width_0_height_0_subtile_0__pin_odata_2_17_,
                   right_width_0_height_0_subtile_0__pin_odata_2_21_,
                   right_width_0_height_0_subtile_0__pin_odata_2_25_,
                   right_width_0_height_0_subtile_0__pin_odata_2_29_,
                   right_width_0_height_0_subtile_0__pin_odata_2_33_,
                   right_width_0_height_0_subtile_0__pin_odata_3_2_,
                   right_width_0_height_0_subtile_0__pin_odata_3_6_,
                   right_width_0_height_0_subtile_0__pin_odata_3_10_,
                   right_width_0_height_0_subtile_0__pin_odata_3_14_,
                   right_width_0_height_0_subtile_0__pin_odata_3_18_,
                   right_width_0_height_0_subtile_0__pin_odata_3_22_,
                   right_width_0_height_0_subtile_0__pin_odata_3_26_,
                   right_width_0_height_0_subtile_0__pin_odata_3_30_,
                   right_width_0_height_0_subtile_0__pin_odata_3_34_,
                   right_width_0_height_0_subtile_0__pin_odata_4_3_,
                   right_width_0_height_0_subtile_0__pin_odata_4_7_,
                   right_width_0_height_0_subtile_0__pin_odata_4_11_,
                   right_width_0_height_0_subtile_0__pin_odata_4_15_,
                   right_width_0_height_0_subtile_0__pin_odata_4_19_,
                   right_width_0_height_0_subtile_0__pin_odata_4_23_,
                   right_width_0_height_0_subtile_0__pin_odata_4_27_,
                   right_width_0_height_0_subtile_0__pin_odata_4_31_,
                   right_width_0_height_0_subtile_0__pin_ovalid_0_0_,
                   right_width_0_height_0_subtile_0__pin_ovalid_4_0_,
                   right_width_0_height_0_subtile_0__pin_ovch_3_0_,
                   right_width_0_height_0_subtile_0__pin_oack_1_0_,
                   right_width_0_height_0_subtile_0__pin_oack_3_0_,
                   right_width_0_height_0_subtile_0__pin_ordy_0_0_,
                   right_width_0_height_0_subtile_0__pin_ordy_2_0_,
                   right_width_0_height_0_subtile_0__pin_ordy_4_0_,
                   right_width_0_height_0_subtile_0__pin_olck_1_0_,
                   right_width_0_height_0_subtile_0__pin_olck_3_0_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_0_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_4_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_8_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_12_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_16_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_20_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_24_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_28_,
                   bottom_width_0_height_0_subtile_0__pin_odata_0_32_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_1_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_5_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_9_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_13_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_17_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_21_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_25_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_29_,
                   bottom_width_0_height_0_subtile_0__pin_odata_1_33_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_2_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_6_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_10_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_14_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_18_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_22_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_26_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_30_,
                   bottom_width_0_height_0_subtile_0__pin_odata_2_34_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_3_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_7_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_11_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_15_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_19_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_23_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_27_,
                   bottom_width_0_height_0_subtile_0__pin_odata_3_31_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_0_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_4_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_8_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_12_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_16_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_20_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_24_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_28_,
                   bottom_width_0_height_0_subtile_0__pin_odata_4_32_,
                   bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_,
                   bottom_width_0_height_0_subtile_0__pin_ovch_0_0_,
                   bottom_width_0_height_0_subtile_0__pin_ovch_4_0_,
                   bottom_width_0_height_0_subtile_0__pin_oack_1_1_,
                   bottom_width_0_height_0_subtile_0__pin_oack_3_1_,
                   bottom_width_0_height_0_subtile_0__pin_ordy_0_1_,
                   bottom_width_0_height_0_subtile_0__pin_ordy_2_1_,
                   bottom_width_0_height_0_subtile_0__pin_ordy_4_1_,
                   bottom_width_0_height_0_subtile_0__pin_olck_1_1_,
                   bottom_width_0_height_0_subtile_0__pin_olck_3_1_,
                   left_width_0_height_0_subtile_0__pin_odata_0_1_,
                   left_width_0_height_0_subtile_0__pin_odata_0_5_,
                   left_width_0_height_0_subtile_0__pin_odata_0_9_,
                   left_width_0_height_0_subtile_0__pin_odata_0_13_,
                   left_width_0_height_0_subtile_0__pin_odata_0_17_,
                   left_width_0_height_0_subtile_0__pin_odata_0_21_,
                   left_width_0_height_0_subtile_0__pin_odata_0_25_,
                   left_width_0_height_0_subtile_0__pin_odata_0_29_,
                   left_width_0_height_0_subtile_0__pin_odata_0_33_,
                   left_width_0_height_0_subtile_0__pin_odata_1_2_,
                   left_width_0_height_0_subtile_0__pin_odata_1_6_,
                   left_width_0_height_0_subtile_0__pin_odata_1_10_,
                   left_width_0_height_0_subtile_0__pin_odata_1_14_,
                   left_width_0_height_0_subtile_0__pin_odata_1_18_,
                   left_width_0_height_0_subtile_0__pin_odata_1_22_,
                   left_width_0_height_0_subtile_0__pin_odata_1_26_,
                   left_width_0_height_0_subtile_0__pin_odata_1_30_,
                   left_width_0_height_0_subtile_0__pin_odata_1_34_,
                   left_width_0_height_0_subtile_0__pin_odata_2_3_,
                   left_width_0_height_0_subtile_0__pin_odata_2_7_,
                   left_width_0_height_0_subtile_0__pin_odata_2_11_,
                   left_width_0_height_0_subtile_0__pin_odata_2_15_,
                   left_width_0_height_0_subtile_0__pin_odata_2_19_,
                   left_width_0_height_0_subtile_0__pin_odata_2_23_,
                   left_width_0_height_0_subtile_0__pin_odata_2_27_,
                   left_width_0_height_0_subtile_0__pin_odata_2_31_,
                   left_width_0_height_0_subtile_0__pin_odata_3_0_,
                   left_width_0_height_0_subtile_0__pin_odata_3_4_,
                   left_width_0_height_0_subtile_0__pin_odata_3_8_,
                   left_width_0_height_0_subtile_0__pin_odata_3_12_,
                   left_width_0_height_0_subtile_0__pin_odata_3_16_,
                   left_width_0_height_0_subtile_0__pin_odata_3_20_,
                   left_width_0_height_0_subtile_0__pin_odata_3_24_,
                   left_width_0_height_0_subtile_0__pin_odata_3_28_,
                   left_width_0_height_0_subtile_0__pin_odata_3_32_,
                   left_width_0_height_0_subtile_0__pin_odata_4_1_,
                   left_width_0_height_0_subtile_0__pin_odata_4_5_,
                   left_width_0_height_0_subtile_0__pin_odata_4_9_,
                   left_width_0_height_0_subtile_0__pin_odata_4_13_,
                   left_width_0_height_0_subtile_0__pin_odata_4_17_,
                   left_width_0_height_0_subtile_0__pin_odata_4_21_,
                   left_width_0_height_0_subtile_0__pin_odata_4_25_,
                   left_width_0_height_0_subtile_0__pin_odata_4_29_,
                   left_width_0_height_0_subtile_0__pin_odata_4_33_,
                   left_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                   left_width_0_height_0_subtile_0__pin_ovch_1_0_,
                   left_width_0_height_0_subtile_0__pin_oack_0_0_,
                   left_width_0_height_0_subtile_0__pin_oack_2_0_,
                   left_width_0_height_0_subtile_0__pin_oack_4_0_,
                   left_width_0_height_0_subtile_0__pin_ordy_1_0_,
                   left_width_0_height_0_subtile_0__pin_ordy_3_0_,
                   left_width_0_height_0_subtile_0__pin_olck_0_0_,
                   left_width_0_height_0_subtile_0__pin_olck_2_0_,
                   left_width_0_height_0_subtile_0__pin_olck_4_0_,
                   ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_rst__0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_my_ypos_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_0_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_4_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_8_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_12_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_16_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_20_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_24_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_28_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_1_32_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_1_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_5_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_9_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_13_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_17_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_21_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_25_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_29_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_2_33_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_2_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_6_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_10_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_14_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_18_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_22_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_26_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_30_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_3_34_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_3_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_7_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_11_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_15_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_19_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_23_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_27_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_idata_4_31_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ivalid_0_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ivalid_4_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ivch_3_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_iack_1_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_iack_3_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ilck_0_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ilck_2_0_;
//----- INPUT PORTS -----
input [0:0] top_width_0_height_0_subtile_0__pin_ilck_4_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_my_xpos_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_20_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_24_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_28_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_0_32_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_5_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_9_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_13_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_17_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_21_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_25_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_29_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_1_33_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_2_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_6_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_10_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_14_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_18_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_22_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_26_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_30_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_2_34_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_3_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_7_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_11_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_15_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_19_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_23_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_27_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_3_31_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_4_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_8_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_12_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_16_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_20_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_24_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_28_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_idata_4_32_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ivalid_1_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ivch_0_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ivch_4_0_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_iack_1_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_iack_3_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ilck_0_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ilck_2_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_ilck_4_1_;
//----- INPUT PORTS -----
input [0:0] right_width_0_height_0_subtile_0__pin_clk_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_my_xpos_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_17_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_21_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_25_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_29_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_0_33_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_2_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_6_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_10_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_14_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_18_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_22_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_26_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_30_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_1_34_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_3_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_7_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_11_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_15_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_19_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_23_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_27_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_2_31_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_4_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_8_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_12_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_16_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_20_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_24_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_28_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_3_32_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_1_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_5_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_9_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_13_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_17_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_21_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_25_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_29_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_idata_4_33_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ivch_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_iack_0_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_iack_2_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_iack_4_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ilck_1_0_;
//----- INPUT PORTS -----
input [0:0] bottom_width_0_height_0_subtile_0__pin_ilck_3_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_my_ypos_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_22_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_26_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_30_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_0_34_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_3_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_7_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_11_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_15_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_19_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_23_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_27_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_1_31_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_4_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_8_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_12_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_16_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_20_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_24_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_28_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_2_32_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_5_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_9_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_13_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_17_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_21_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_25_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_29_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_3_33_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_2_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_6_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_10_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_14_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_18_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_22_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_26_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_30_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_idata_4_34_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_ivalid_3_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_ivch_2_0_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_iack_0_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_iack_2_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_iack_4_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_ilck_1_1_;
//----- INPUT PORTS -----
input [0:0] left_width_0_height_0_subtile_0__pin_ilck_3_1_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_14_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_18_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_22_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_26_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_30_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_0_34_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_3_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_7_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_11_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_15_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_19_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_23_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_27_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_1_31_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_4_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_8_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_12_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_16_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_20_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_24_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_28_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_2_32_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_5_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_9_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_13_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_17_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_21_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_25_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_29_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_3_33_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_2_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_6_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_10_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_14_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_18_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_22_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_26_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_30_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_odata_4_34_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_ovalid_3_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_ovch_2_0_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_oack_0_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_oack_2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_oack_4_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_ordy_1_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_ordy_3_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_olck_0_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_olck_2_1_;
//----- OUTPUT PORTS -----
output [0:0] top_width_0_height_0_subtile_0__pin_olck_4_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_27_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_0_31_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_4_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_8_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_12_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_16_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_20_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_24_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_28_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_1_32_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_1_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_5_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_9_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_13_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_17_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_21_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_25_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_29_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_2_33_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_2_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_6_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_10_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_14_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_18_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_22_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_26_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_30_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_3_34_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_3_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_7_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_11_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_15_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_19_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_23_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_27_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_odata_4_31_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ovalid_0_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ovalid_4_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ovch_3_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_oack_1_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_oack_3_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ordy_0_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ordy_2_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_ordy_4_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_olck_1_0_;
//----- OUTPUT PORTS -----
output [0:0] right_width_0_height_0_subtile_0__pin_olck_3_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
//----- OUTPUT PORTS -----
output [0:0] bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_9_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_13_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_17_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_21_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_25_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_29_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_0_33_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_2_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_6_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_10_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_14_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_18_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_22_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_26_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_30_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_1_34_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_4_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_8_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_12_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_16_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_20_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_24_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_28_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_3_32_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_1_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_5_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_9_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_13_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_17_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_21_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_25_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_29_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_odata_4_33_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_ovch_1_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_oack_0_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_oack_4_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_ordy_1_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_ordy_3_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_olck_0_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- OUTPUT PORTS -----
output [0:0] left_width_0_height_0_subtile_0__pin_olck_4_0_;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----



// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_router_mode_router_ logical_tile_router_mode_router__0 (
		.clk(clk),
		.set(set),
		.reset(reset),
		.prog_clk(prog_clk),
		.router_rst_(top_width_0_height_0_subtile_0__pin_rst__0_),
		.router_my_xpos({right_width_0_height_0_subtile_0__pin_my_xpos_0_, bottom_width_0_height_0_subtile_0__pin_my_xpos_1_}),
		.router_my_ypos({left_width_0_height_0_subtile_0__pin_my_ypos_0_, top_width_0_height_0_subtile_0__pin_my_ypos_1_}),
		.router_idata_0({right_width_0_height_0_subtile_0__pin_idata_0_0_, bottom_width_0_height_0_subtile_0__pin_idata_0_1_, left_width_0_height_0_subtile_0__pin_idata_0_2_, top_width_0_height_0_subtile_0__pin_idata_0_3_, right_width_0_height_0_subtile_0__pin_idata_0_4_, bottom_width_0_height_0_subtile_0__pin_idata_0_5_, left_width_0_height_0_subtile_0__pin_idata_0_6_, top_width_0_height_0_subtile_0__pin_idata_0_7_, right_width_0_height_0_subtile_0__pin_idata_0_8_, bottom_width_0_height_0_subtile_0__pin_idata_0_9_, left_width_0_height_0_subtile_0__pin_idata_0_10_, top_width_0_height_0_subtile_0__pin_idata_0_11_, right_width_0_height_0_subtile_0__pin_idata_0_12_, bottom_width_0_height_0_subtile_0__pin_idata_0_13_, left_width_0_height_0_subtile_0__pin_idata_0_14_, top_width_0_height_0_subtile_0__pin_idata_0_15_, right_width_0_height_0_subtile_0__pin_idata_0_16_, bottom_width_0_height_0_subtile_0__pin_idata_0_17_, left_width_0_height_0_subtile_0__pin_idata_0_18_, top_width_0_height_0_subtile_0__pin_idata_0_19_, right_width_0_height_0_subtile_0__pin_idata_0_20_, bottom_width_0_height_0_subtile_0__pin_idata_0_21_, left_width_0_height_0_subtile_0__pin_idata_0_22_, top_width_0_height_0_subtile_0__pin_idata_0_23_, right_width_0_height_0_subtile_0__pin_idata_0_24_, bottom_width_0_height_0_subtile_0__pin_idata_0_25_, left_width_0_height_0_subtile_0__pin_idata_0_26_, top_width_0_height_0_subtile_0__pin_idata_0_27_, right_width_0_height_0_subtile_0__pin_idata_0_28_, bottom_width_0_height_0_subtile_0__pin_idata_0_29_, left_width_0_height_0_subtile_0__pin_idata_0_30_, top_width_0_height_0_subtile_0__pin_idata_0_31_, right_width_0_height_0_subtile_0__pin_idata_0_32_, bottom_width_0_height_0_subtile_0__pin_idata_0_33_, left_width_0_height_0_subtile_0__pin_idata_0_34_}),
		.router_idata_1({top_width_0_height_0_subtile_0__pin_idata_1_0_, right_width_0_height_0_subtile_0__pin_idata_1_1_, bottom_width_0_height_0_subtile_0__pin_idata_1_2_, left_width_0_height_0_subtile_0__pin_idata_1_3_, top_width_0_height_0_subtile_0__pin_idata_1_4_, right_width_0_height_0_subtile_0__pin_idata_1_5_, bottom_width_0_height_0_subtile_0__pin_idata_1_6_, left_width_0_height_0_subtile_0__pin_idata_1_7_, top_width_0_height_0_subtile_0__pin_idata_1_8_, right_width_0_height_0_subtile_0__pin_idata_1_9_, bottom_width_0_height_0_subtile_0__pin_idata_1_10_, left_width_0_height_0_subtile_0__pin_idata_1_11_, top_width_0_height_0_subtile_0__pin_idata_1_12_, right_width_0_height_0_subtile_0__pin_idata_1_13_, bottom_width_0_height_0_subtile_0__pin_idata_1_14_, left_width_0_height_0_subtile_0__pin_idata_1_15_, top_width_0_height_0_subtile_0__pin_idata_1_16_, right_width_0_height_0_subtile_0__pin_idata_1_17_, bottom_width_0_height_0_subtile_0__pin_idata_1_18_, left_width_0_height_0_subtile_0__pin_idata_1_19_, top_width_0_height_0_subtile_0__pin_idata_1_20_, right_width_0_height_0_subtile_0__pin_idata_1_21_, bottom_width_0_height_0_subtile_0__pin_idata_1_22_, left_width_0_height_0_subtile_0__pin_idata_1_23_, top_width_0_height_0_subtile_0__pin_idata_1_24_, right_width_0_height_0_subtile_0__pin_idata_1_25_, bottom_width_0_height_0_subtile_0__pin_idata_1_26_, left_width_0_height_0_subtile_0__pin_idata_1_27_, top_width_0_height_0_subtile_0__pin_idata_1_28_, right_width_0_height_0_subtile_0__pin_idata_1_29_, bottom_width_0_height_0_subtile_0__pin_idata_1_30_, left_width_0_height_0_subtile_0__pin_idata_1_31_, top_width_0_height_0_subtile_0__pin_idata_1_32_, right_width_0_height_0_subtile_0__pin_idata_1_33_, bottom_width_0_height_0_subtile_0__pin_idata_1_34_}),
		.router_idata_2({left_width_0_height_0_subtile_0__pin_idata_2_0_, top_width_0_height_0_subtile_0__pin_idata_2_1_, right_width_0_height_0_subtile_0__pin_idata_2_2_, bottom_width_0_height_0_subtile_0__pin_idata_2_3_, left_width_0_height_0_subtile_0__pin_idata_2_4_, top_width_0_height_0_subtile_0__pin_idata_2_5_, right_width_0_height_0_subtile_0__pin_idata_2_6_, bottom_width_0_height_0_subtile_0__pin_idata_2_7_, left_width_0_height_0_subtile_0__pin_idata_2_8_, top_width_0_height_0_subtile_0__pin_idata_2_9_, right_width_0_height_0_subtile_0__pin_idata_2_10_, bottom_width_0_height_0_subtile_0__pin_idata_2_11_, left_width_0_height_0_subtile_0__pin_idata_2_12_, top_width_0_height_0_subtile_0__pin_idata_2_13_, right_width_0_height_0_subtile_0__pin_idata_2_14_, bottom_width_0_height_0_subtile_0__pin_idata_2_15_, left_width_0_height_0_subtile_0__pin_idata_2_16_, top_width_0_height_0_subtile_0__pin_idata_2_17_, right_width_0_height_0_subtile_0__pin_idata_2_18_, bottom_width_0_height_0_subtile_0__pin_idata_2_19_, left_width_0_height_0_subtile_0__pin_idata_2_20_, top_width_0_height_0_subtile_0__pin_idata_2_21_, right_width_0_height_0_subtile_0__pin_idata_2_22_, bottom_width_0_height_0_subtile_0__pin_idata_2_23_, left_width_0_height_0_subtile_0__pin_idata_2_24_, top_width_0_height_0_subtile_0__pin_idata_2_25_, right_width_0_height_0_subtile_0__pin_idata_2_26_, bottom_width_0_height_0_subtile_0__pin_idata_2_27_, left_width_0_height_0_subtile_0__pin_idata_2_28_, top_width_0_height_0_subtile_0__pin_idata_2_29_, right_width_0_height_0_subtile_0__pin_idata_2_30_, bottom_width_0_height_0_subtile_0__pin_idata_2_31_, left_width_0_height_0_subtile_0__pin_idata_2_32_, top_width_0_height_0_subtile_0__pin_idata_2_33_, right_width_0_height_0_subtile_0__pin_idata_2_34_}),
		.router_idata_3({bottom_width_0_height_0_subtile_0__pin_idata_3_0_, left_width_0_height_0_subtile_0__pin_idata_3_1_, top_width_0_height_0_subtile_0__pin_idata_3_2_, right_width_0_height_0_subtile_0__pin_idata_3_3_, bottom_width_0_height_0_subtile_0__pin_idata_3_4_, left_width_0_height_0_subtile_0__pin_idata_3_5_, top_width_0_height_0_subtile_0__pin_idata_3_6_, right_width_0_height_0_subtile_0__pin_idata_3_7_, bottom_width_0_height_0_subtile_0__pin_idata_3_8_, left_width_0_height_0_subtile_0__pin_idata_3_9_, top_width_0_height_0_subtile_0__pin_idata_3_10_, right_width_0_height_0_subtile_0__pin_idata_3_11_, bottom_width_0_height_0_subtile_0__pin_idata_3_12_, left_width_0_height_0_subtile_0__pin_idata_3_13_, top_width_0_height_0_subtile_0__pin_idata_3_14_, right_width_0_height_0_subtile_0__pin_idata_3_15_, bottom_width_0_height_0_subtile_0__pin_idata_3_16_, left_width_0_height_0_subtile_0__pin_idata_3_17_, top_width_0_height_0_subtile_0__pin_idata_3_18_, right_width_0_height_0_subtile_0__pin_idata_3_19_, bottom_width_0_height_0_subtile_0__pin_idata_3_20_, left_width_0_height_0_subtile_0__pin_idata_3_21_, top_width_0_height_0_subtile_0__pin_idata_3_22_, right_width_0_height_0_subtile_0__pin_idata_3_23_, bottom_width_0_height_0_subtile_0__pin_idata_3_24_, left_width_0_height_0_subtile_0__pin_idata_3_25_, top_width_0_height_0_subtile_0__pin_idata_3_26_, right_width_0_height_0_subtile_0__pin_idata_3_27_, bottom_width_0_height_0_subtile_0__pin_idata_3_28_, left_width_0_height_0_subtile_0__pin_idata_3_29_, top_width_0_height_0_subtile_0__pin_idata_3_30_, right_width_0_height_0_subtile_0__pin_idata_3_31_, bottom_width_0_height_0_subtile_0__pin_idata_3_32_, left_width_0_height_0_subtile_0__pin_idata_3_33_, top_width_0_height_0_subtile_0__pin_idata_3_34_}),
		.router_idata_4({right_width_0_height_0_subtile_0__pin_idata_4_0_, bottom_width_0_height_0_subtile_0__pin_idata_4_1_, left_width_0_height_0_subtile_0__pin_idata_4_2_, top_width_0_height_0_subtile_0__pin_idata_4_3_, right_width_0_height_0_subtile_0__pin_idata_4_4_, bottom_width_0_height_0_subtile_0__pin_idata_4_5_, left_width_0_height_0_subtile_0__pin_idata_4_6_, top_width_0_height_0_subtile_0__pin_idata_4_7_, right_width_0_height_0_subtile_0__pin_idata_4_8_, bottom_width_0_height_0_subtile_0__pin_idata_4_9_, left_width_0_height_0_subtile_0__pin_idata_4_10_, top_width_0_height_0_subtile_0__pin_idata_4_11_, right_width_0_height_0_subtile_0__pin_idata_4_12_, bottom_width_0_height_0_subtile_0__pin_idata_4_13_, left_width_0_height_0_subtile_0__pin_idata_4_14_, top_width_0_height_0_subtile_0__pin_idata_4_15_, right_width_0_height_0_subtile_0__pin_idata_4_16_, bottom_width_0_height_0_subtile_0__pin_idata_4_17_, left_width_0_height_0_subtile_0__pin_idata_4_18_, top_width_0_height_0_subtile_0__pin_idata_4_19_, right_width_0_height_0_subtile_0__pin_idata_4_20_, bottom_width_0_height_0_subtile_0__pin_idata_4_21_, left_width_0_height_0_subtile_0__pin_idata_4_22_, top_width_0_height_0_subtile_0__pin_idata_4_23_, right_width_0_height_0_subtile_0__pin_idata_4_24_, bottom_width_0_height_0_subtile_0__pin_idata_4_25_, left_width_0_height_0_subtile_0__pin_idata_4_26_, top_width_0_height_0_subtile_0__pin_idata_4_27_, right_width_0_height_0_subtile_0__pin_idata_4_28_, bottom_width_0_height_0_subtile_0__pin_idata_4_29_, left_width_0_height_0_subtile_0__pin_idata_4_30_, top_width_0_height_0_subtile_0__pin_idata_4_31_, right_width_0_height_0_subtile_0__pin_idata_4_32_, bottom_width_0_height_0_subtile_0__pin_idata_4_33_, left_width_0_height_0_subtile_0__pin_idata_4_34_}),
		.router_ivalid_0(top_width_0_height_0_subtile_0__pin_ivalid_0_0_),
		.router_ivalid_1(right_width_0_height_0_subtile_0__pin_ivalid_1_0_),
		.router_ivalid_2(bottom_width_0_height_0_subtile_0__pin_ivalid_2_0_),
		.router_ivalid_3(left_width_0_height_0_subtile_0__pin_ivalid_3_0_),
		.router_ivalid_4(top_width_0_height_0_subtile_0__pin_ivalid_4_0_),
		.router_ivch_0(right_width_0_height_0_subtile_0__pin_ivch_0_0_),
		.router_ivch_1(bottom_width_0_height_0_subtile_0__pin_ivch_1_0_),
		.router_ivch_2(left_width_0_height_0_subtile_0__pin_ivch_2_0_),
		.router_ivch_3(top_width_0_height_0_subtile_0__pin_ivch_3_0_),
		.router_ivch_4(right_width_0_height_0_subtile_0__pin_ivch_4_0_),
		.router_iack_0({bottom_width_0_height_0_subtile_0__pin_iack_0_0_, left_width_0_height_0_subtile_0__pin_iack_0_1_}),
		.router_iack_1({top_width_0_height_0_subtile_0__pin_iack_1_0_, right_width_0_height_0_subtile_0__pin_iack_1_1_}),
		.router_iack_2({bottom_width_0_height_0_subtile_0__pin_iack_2_0_, left_width_0_height_0_subtile_0__pin_iack_2_1_}),
		.router_iack_3({top_width_0_height_0_subtile_0__pin_iack_3_0_, right_width_0_height_0_subtile_0__pin_iack_3_1_}),
		.router_iack_4({bottom_width_0_height_0_subtile_0__pin_iack_4_0_, left_width_0_height_0_subtile_0__pin_iack_4_1_}),
		.router_ilck_0({top_width_0_height_0_subtile_0__pin_ilck_0_0_, right_width_0_height_0_subtile_0__pin_ilck_0_1_}),
		.router_ilck_1({bottom_width_0_height_0_subtile_0__pin_ilck_1_0_, left_width_0_height_0_subtile_0__pin_ilck_1_1_}),
		.router_ilck_2({top_width_0_height_0_subtile_0__pin_ilck_2_0_, right_width_0_height_0_subtile_0__pin_ilck_2_1_}),
		.router_ilck_3({bottom_width_0_height_0_subtile_0__pin_ilck_3_0_, left_width_0_height_0_subtile_0__pin_ilck_3_1_}),
		.router_ilck_4({top_width_0_height_0_subtile_0__pin_ilck_4_0_, right_width_0_height_0_subtile_0__pin_ilck_4_1_}),
		.router_clk(right_width_0_height_0_subtile_0__pin_clk_0_),
		.ccff_head(ccff_head),
		.router_odata_0({bottom_width_0_height_0_subtile_0__pin_odata_0_0_, left_width_0_height_0_subtile_0__pin_odata_0_1_, top_width_0_height_0_subtile_0__pin_odata_0_2_, right_width_0_height_0_subtile_0__pin_odata_0_3_, bottom_width_0_height_0_subtile_0__pin_odata_0_4_, left_width_0_height_0_subtile_0__pin_odata_0_5_, top_width_0_height_0_subtile_0__pin_odata_0_6_, right_width_0_height_0_subtile_0__pin_odata_0_7_, bottom_width_0_height_0_subtile_0__pin_odata_0_8_, left_width_0_height_0_subtile_0__pin_odata_0_9_, top_width_0_height_0_subtile_0__pin_odata_0_10_, right_width_0_height_0_subtile_0__pin_odata_0_11_, bottom_width_0_height_0_subtile_0__pin_odata_0_12_, left_width_0_height_0_subtile_0__pin_odata_0_13_, top_width_0_height_0_subtile_0__pin_odata_0_14_, right_width_0_height_0_subtile_0__pin_odata_0_15_, bottom_width_0_height_0_subtile_0__pin_odata_0_16_, left_width_0_height_0_subtile_0__pin_odata_0_17_, top_width_0_height_0_subtile_0__pin_odata_0_18_, right_width_0_height_0_subtile_0__pin_odata_0_19_, bottom_width_0_height_0_subtile_0__pin_odata_0_20_, left_width_0_height_0_subtile_0__pin_odata_0_21_, top_width_0_height_0_subtile_0__pin_odata_0_22_, right_width_0_height_0_subtile_0__pin_odata_0_23_, bottom_width_0_height_0_subtile_0__pin_odata_0_24_, left_width_0_height_0_subtile_0__pin_odata_0_25_, top_width_0_height_0_subtile_0__pin_odata_0_26_, right_width_0_height_0_subtile_0__pin_odata_0_27_, bottom_width_0_height_0_subtile_0__pin_odata_0_28_, left_width_0_height_0_subtile_0__pin_odata_0_29_, top_width_0_height_0_subtile_0__pin_odata_0_30_, right_width_0_height_0_subtile_0__pin_odata_0_31_, bottom_width_0_height_0_subtile_0__pin_odata_0_32_, left_width_0_height_0_subtile_0__pin_odata_0_33_, top_width_0_height_0_subtile_0__pin_odata_0_34_}),
		.router_odata_1({right_width_0_height_0_subtile_0__pin_odata_1_0_, bottom_width_0_height_0_subtile_0__pin_odata_1_1_, left_width_0_height_0_subtile_0__pin_odata_1_2_, top_width_0_height_0_subtile_0__pin_odata_1_3_, right_width_0_height_0_subtile_0__pin_odata_1_4_, bottom_width_0_height_0_subtile_0__pin_odata_1_5_, left_width_0_height_0_subtile_0__pin_odata_1_6_, top_width_0_height_0_subtile_0__pin_odata_1_7_, right_width_0_height_0_subtile_0__pin_odata_1_8_, bottom_width_0_height_0_subtile_0__pin_odata_1_9_, left_width_0_height_0_subtile_0__pin_odata_1_10_, top_width_0_height_0_subtile_0__pin_odata_1_11_, right_width_0_height_0_subtile_0__pin_odata_1_12_, bottom_width_0_height_0_subtile_0__pin_odata_1_13_, left_width_0_height_0_subtile_0__pin_odata_1_14_, top_width_0_height_0_subtile_0__pin_odata_1_15_, right_width_0_height_0_subtile_0__pin_odata_1_16_, bottom_width_0_height_0_subtile_0__pin_odata_1_17_, left_width_0_height_0_subtile_0__pin_odata_1_18_, top_width_0_height_0_subtile_0__pin_odata_1_19_, right_width_0_height_0_subtile_0__pin_odata_1_20_, bottom_width_0_height_0_subtile_0__pin_odata_1_21_, left_width_0_height_0_subtile_0__pin_odata_1_22_, top_width_0_height_0_subtile_0__pin_odata_1_23_, right_width_0_height_0_subtile_0__pin_odata_1_24_, bottom_width_0_height_0_subtile_0__pin_odata_1_25_, left_width_0_height_0_subtile_0__pin_odata_1_26_, top_width_0_height_0_subtile_0__pin_odata_1_27_, right_width_0_height_0_subtile_0__pin_odata_1_28_, bottom_width_0_height_0_subtile_0__pin_odata_1_29_, left_width_0_height_0_subtile_0__pin_odata_1_30_, top_width_0_height_0_subtile_0__pin_odata_1_31_, right_width_0_height_0_subtile_0__pin_odata_1_32_, bottom_width_0_height_0_subtile_0__pin_odata_1_33_, left_width_0_height_0_subtile_0__pin_odata_1_34_}),
		.router_odata_2({top_width_0_height_0_subtile_0__pin_odata_2_0_, right_width_0_height_0_subtile_0__pin_odata_2_1_, bottom_width_0_height_0_subtile_0__pin_odata_2_2_, left_width_0_height_0_subtile_0__pin_odata_2_3_, top_width_0_height_0_subtile_0__pin_odata_2_4_, right_width_0_height_0_subtile_0__pin_odata_2_5_, bottom_width_0_height_0_subtile_0__pin_odata_2_6_, left_width_0_height_0_subtile_0__pin_odata_2_7_, top_width_0_height_0_subtile_0__pin_odata_2_8_, right_width_0_height_0_subtile_0__pin_odata_2_9_, bottom_width_0_height_0_subtile_0__pin_odata_2_10_, left_width_0_height_0_subtile_0__pin_odata_2_11_, top_width_0_height_0_subtile_0__pin_odata_2_12_, right_width_0_height_0_subtile_0__pin_odata_2_13_, bottom_width_0_height_0_subtile_0__pin_odata_2_14_, left_width_0_height_0_subtile_0__pin_odata_2_15_, top_width_0_height_0_subtile_0__pin_odata_2_16_, right_width_0_height_0_subtile_0__pin_odata_2_17_, bottom_width_0_height_0_subtile_0__pin_odata_2_18_, left_width_0_height_0_subtile_0__pin_odata_2_19_, top_width_0_height_0_subtile_0__pin_odata_2_20_, right_width_0_height_0_subtile_0__pin_odata_2_21_, bottom_width_0_height_0_subtile_0__pin_odata_2_22_, left_width_0_height_0_subtile_0__pin_odata_2_23_, top_width_0_height_0_subtile_0__pin_odata_2_24_, right_width_0_height_0_subtile_0__pin_odata_2_25_, bottom_width_0_height_0_subtile_0__pin_odata_2_26_, left_width_0_height_0_subtile_0__pin_odata_2_27_, top_width_0_height_0_subtile_0__pin_odata_2_28_, right_width_0_height_0_subtile_0__pin_odata_2_29_, bottom_width_0_height_0_subtile_0__pin_odata_2_30_, left_width_0_height_0_subtile_0__pin_odata_2_31_, top_width_0_height_0_subtile_0__pin_odata_2_32_, right_width_0_height_0_subtile_0__pin_odata_2_33_, bottom_width_0_height_0_subtile_0__pin_odata_2_34_}),
		.router_odata_3({left_width_0_height_0_subtile_0__pin_odata_3_0_, top_width_0_height_0_subtile_0__pin_odata_3_1_, right_width_0_height_0_subtile_0__pin_odata_3_2_, bottom_width_0_height_0_subtile_0__pin_odata_3_3_, left_width_0_height_0_subtile_0__pin_odata_3_4_, top_width_0_height_0_subtile_0__pin_odata_3_5_, right_width_0_height_0_subtile_0__pin_odata_3_6_, bottom_width_0_height_0_subtile_0__pin_odata_3_7_, left_width_0_height_0_subtile_0__pin_odata_3_8_, top_width_0_height_0_subtile_0__pin_odata_3_9_, right_width_0_height_0_subtile_0__pin_odata_3_10_, bottom_width_0_height_0_subtile_0__pin_odata_3_11_, left_width_0_height_0_subtile_0__pin_odata_3_12_, top_width_0_height_0_subtile_0__pin_odata_3_13_, right_width_0_height_0_subtile_0__pin_odata_3_14_, bottom_width_0_height_0_subtile_0__pin_odata_3_15_, left_width_0_height_0_subtile_0__pin_odata_3_16_, top_width_0_height_0_subtile_0__pin_odata_3_17_, right_width_0_height_0_subtile_0__pin_odata_3_18_, bottom_width_0_height_0_subtile_0__pin_odata_3_19_, left_width_0_height_0_subtile_0__pin_odata_3_20_, top_width_0_height_0_subtile_0__pin_odata_3_21_, right_width_0_height_0_subtile_0__pin_odata_3_22_, bottom_width_0_height_0_subtile_0__pin_odata_3_23_, left_width_0_height_0_subtile_0__pin_odata_3_24_, top_width_0_height_0_subtile_0__pin_odata_3_25_, right_width_0_height_0_subtile_0__pin_odata_3_26_, bottom_width_0_height_0_subtile_0__pin_odata_3_27_, left_width_0_height_0_subtile_0__pin_odata_3_28_, top_width_0_height_0_subtile_0__pin_odata_3_29_, right_width_0_height_0_subtile_0__pin_odata_3_30_, bottom_width_0_height_0_subtile_0__pin_odata_3_31_, left_width_0_height_0_subtile_0__pin_odata_3_32_, top_width_0_height_0_subtile_0__pin_odata_3_33_, right_width_0_height_0_subtile_0__pin_odata_3_34_}),
		.router_odata_4({bottom_width_0_height_0_subtile_0__pin_odata_4_0_, left_width_0_height_0_subtile_0__pin_odata_4_1_, top_width_0_height_0_subtile_0__pin_odata_4_2_, right_width_0_height_0_subtile_0__pin_odata_4_3_, bottom_width_0_height_0_subtile_0__pin_odata_4_4_, left_width_0_height_0_subtile_0__pin_odata_4_5_, top_width_0_height_0_subtile_0__pin_odata_4_6_, right_width_0_height_0_subtile_0__pin_odata_4_7_, bottom_width_0_height_0_subtile_0__pin_odata_4_8_, left_width_0_height_0_subtile_0__pin_odata_4_9_, top_width_0_height_0_subtile_0__pin_odata_4_10_, right_width_0_height_0_subtile_0__pin_odata_4_11_, bottom_width_0_height_0_subtile_0__pin_odata_4_12_, left_width_0_height_0_subtile_0__pin_odata_4_13_, top_width_0_height_0_subtile_0__pin_odata_4_14_, right_width_0_height_0_subtile_0__pin_odata_4_15_, bottom_width_0_height_0_subtile_0__pin_odata_4_16_, left_width_0_height_0_subtile_0__pin_odata_4_17_, top_width_0_height_0_subtile_0__pin_odata_4_18_, right_width_0_height_0_subtile_0__pin_odata_4_19_, bottom_width_0_height_0_subtile_0__pin_odata_4_20_, left_width_0_height_0_subtile_0__pin_odata_4_21_, top_width_0_height_0_subtile_0__pin_odata_4_22_, right_width_0_height_0_subtile_0__pin_odata_4_23_, bottom_width_0_height_0_subtile_0__pin_odata_4_24_, left_width_0_height_0_subtile_0__pin_odata_4_25_, top_width_0_height_0_subtile_0__pin_odata_4_26_, right_width_0_height_0_subtile_0__pin_odata_4_27_, bottom_width_0_height_0_subtile_0__pin_odata_4_28_, left_width_0_height_0_subtile_0__pin_odata_4_29_, top_width_0_height_0_subtile_0__pin_odata_4_30_, right_width_0_height_0_subtile_0__pin_odata_4_31_, bottom_width_0_height_0_subtile_0__pin_odata_4_32_, left_width_0_height_0_subtile_0__pin_odata_4_33_, top_width_0_height_0_subtile_0__pin_odata_4_34_}),
		.router_ovalid_0(right_width_0_height_0_subtile_0__pin_ovalid_0_0_),
		.router_ovalid_1(bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_),
		.router_ovalid_2(left_width_0_height_0_subtile_0__pin_ovalid_2_0_),
		.router_ovalid_3(top_width_0_height_0_subtile_0__pin_ovalid_3_0_),
		.router_ovalid_4(right_width_0_height_0_subtile_0__pin_ovalid_4_0_),
		.router_ovch_0(bottom_width_0_height_0_subtile_0__pin_ovch_0_0_),
		.router_ovch_1(left_width_0_height_0_subtile_0__pin_ovch_1_0_),
		.router_ovch_2(top_width_0_height_0_subtile_0__pin_ovch_2_0_),
		.router_ovch_3(right_width_0_height_0_subtile_0__pin_ovch_3_0_),
		.router_ovch_4(bottom_width_0_height_0_subtile_0__pin_ovch_4_0_),
		.router_oack_0({left_width_0_height_0_subtile_0__pin_oack_0_0_, top_width_0_height_0_subtile_0__pin_oack_0_1_}),
		.router_oack_1({right_width_0_height_0_subtile_0__pin_oack_1_0_, bottom_width_0_height_0_subtile_0__pin_oack_1_1_}),
		.router_oack_2({left_width_0_height_0_subtile_0__pin_oack_2_0_, top_width_0_height_0_subtile_0__pin_oack_2_1_}),
		.router_oack_3({right_width_0_height_0_subtile_0__pin_oack_3_0_, bottom_width_0_height_0_subtile_0__pin_oack_3_1_}),
		.router_oack_4({left_width_0_height_0_subtile_0__pin_oack_4_0_, top_width_0_height_0_subtile_0__pin_oack_4_1_}),
		.router_ordy_0({right_width_0_height_0_subtile_0__pin_ordy_0_0_, bottom_width_0_height_0_subtile_0__pin_ordy_0_1_}),
		.router_ordy_1({left_width_0_height_0_subtile_0__pin_ordy_1_0_, top_width_0_height_0_subtile_0__pin_ordy_1_1_}),
		.router_ordy_2({right_width_0_height_0_subtile_0__pin_ordy_2_0_, bottom_width_0_height_0_subtile_0__pin_ordy_2_1_}),
		.router_ordy_3({left_width_0_height_0_subtile_0__pin_ordy_3_0_, top_width_0_height_0_subtile_0__pin_ordy_3_1_}),
		.router_ordy_4({right_width_0_height_0_subtile_0__pin_ordy_4_0_, bottom_width_0_height_0_subtile_0__pin_ordy_4_1_}),
		.router_olck_0({left_width_0_height_0_subtile_0__pin_olck_0_0_, top_width_0_height_0_subtile_0__pin_olck_0_1_}),
		.router_olck_1({right_width_0_height_0_subtile_0__pin_olck_1_0_, bottom_width_0_height_0_subtile_0__pin_olck_1_1_}),
		.router_olck_2({left_width_0_height_0_subtile_0__pin_olck_2_0_, top_width_0_height_0_subtile_0__pin_olck_2_1_}),
		.router_olck_3({right_width_0_height_0_subtile_0__pin_olck_3_0_, bottom_width_0_height_0_subtile_0__pin_olck_3_1_}),
		.router_olck_4({left_width_0_height_0_subtile_0__pin_olck_4_0_, top_width_0_height_0_subtile_0__pin_olck_4_1_}),
		.ccff_tail(ccff_tail));

endmodule
// ----- END Verilog module for grid_router -----

//----- Default net type -----
`default_nettype wire



// ----- END Grid Verilog module: grid_router -----

