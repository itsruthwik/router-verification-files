//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[5][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jul  5 01:26:08 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_5__5_ -----
module sb_5__5_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:284] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_;
//----- INPUT PORTS -----
input [0:284] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:284] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:284] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:284] chany_top_out;
//----- OUTPUT PORTS -----
output [0:284] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:284] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:284] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size15_0_sram;
wire [0:3] mux_tree_tapbuf_size15_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_1_sram;
wire [0:3] mux_tree_tapbuf_size15_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_1_ccff_tail;
wire [0:4] mux_tree_tapbuf_size16_0_sram;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_10_sram;
wire [0:4] mux_tree_tapbuf_size16_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_11_sram;
wire [0:4] mux_tree_tapbuf_size16_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_12_sram;
wire [0:4] mux_tree_tapbuf_size16_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_13_sram;
wire [0:4] mux_tree_tapbuf_size16_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_14_sram;
wire [0:4] mux_tree_tapbuf_size16_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_15_sram;
wire [0:4] mux_tree_tapbuf_size16_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_16_sram;
wire [0:4] mux_tree_tapbuf_size16_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_17_sram;
wire [0:4] mux_tree_tapbuf_size16_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_18_sram;
wire [0:4] mux_tree_tapbuf_size16_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_19_sram;
wire [0:4] mux_tree_tapbuf_size16_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_1_sram;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_20_sram;
wire [0:4] mux_tree_tapbuf_size16_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_21_sram;
wire [0:4] mux_tree_tapbuf_size16_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_22_sram;
wire [0:4] mux_tree_tapbuf_size16_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_23_sram;
wire [0:4] mux_tree_tapbuf_size16_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_24_sram;
wire [0:4] mux_tree_tapbuf_size16_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_25_sram;
wire [0:4] mux_tree_tapbuf_size16_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_26_sram;
wire [0:4] mux_tree_tapbuf_size16_26_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_27_sram;
wire [0:4] mux_tree_tapbuf_size16_27_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_28_sram;
wire [0:4] mux_tree_tapbuf_size16_28_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_29_sram;
wire [0:4] mux_tree_tapbuf_size16_29_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_2_sram;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_30_sram;
wire [0:4] mux_tree_tapbuf_size16_30_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_31_sram;
wire [0:4] mux_tree_tapbuf_size16_31_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_32_sram;
wire [0:4] mux_tree_tapbuf_size16_32_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_33_sram;
wire [0:4] mux_tree_tapbuf_size16_33_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_34_sram;
wire [0:4] mux_tree_tapbuf_size16_34_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_35_sram;
wire [0:4] mux_tree_tapbuf_size16_35_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_36_sram;
wire [0:4] mux_tree_tapbuf_size16_36_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_37_sram;
wire [0:4] mux_tree_tapbuf_size16_37_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_38_sram;
wire [0:4] mux_tree_tapbuf_size16_38_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_39_sram;
wire [0:4] mux_tree_tapbuf_size16_39_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_3_sram;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_40_sram;
wire [0:4] mux_tree_tapbuf_size16_40_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_41_sram;
wire [0:4] mux_tree_tapbuf_size16_41_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_42_sram;
wire [0:4] mux_tree_tapbuf_size16_42_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_43_sram;
wire [0:4] mux_tree_tapbuf_size16_43_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_44_sram;
wire [0:4] mux_tree_tapbuf_size16_44_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_45_sram;
wire [0:4] mux_tree_tapbuf_size16_45_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_46_sram;
wire [0:4] mux_tree_tapbuf_size16_46_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_4_sram;
wire [0:4] mux_tree_tapbuf_size16_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_5_sram;
wire [0:4] mux_tree_tapbuf_size16_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_6_sram;
wire [0:4] mux_tree_tapbuf_size16_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_7_sram;
wire [0:4] mux_tree_tapbuf_size16_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_8_sram;
wire [0:4] mux_tree_tapbuf_size16_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_9_sram;
wire [0:4] mux_tree_tapbuf_size16_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size17_0_sram;
wire [0:4] mux_tree_tapbuf_size17_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_10_sram;
wire [0:4] mux_tree_tapbuf_size17_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_11_sram;
wire [0:4] mux_tree_tapbuf_size17_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_12_sram;
wire [0:4] mux_tree_tapbuf_size17_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_13_sram;
wire [0:4] mux_tree_tapbuf_size17_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_14_sram;
wire [0:4] mux_tree_tapbuf_size17_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_15_sram;
wire [0:4] mux_tree_tapbuf_size17_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_16_sram;
wire [0:4] mux_tree_tapbuf_size17_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_17_sram;
wire [0:4] mux_tree_tapbuf_size17_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_18_sram;
wire [0:4] mux_tree_tapbuf_size17_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_19_sram;
wire [0:4] mux_tree_tapbuf_size17_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_1_sram;
wire [0:4] mux_tree_tapbuf_size17_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_20_sram;
wire [0:4] mux_tree_tapbuf_size17_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_21_sram;
wire [0:4] mux_tree_tapbuf_size17_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_2_sram;
wire [0:4] mux_tree_tapbuf_size17_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_3_sram;
wire [0:4] mux_tree_tapbuf_size17_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_4_sram;
wire [0:4] mux_tree_tapbuf_size17_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_5_sram;
wire [0:4] mux_tree_tapbuf_size17_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_6_sram;
wire [0:4] mux_tree_tapbuf_size17_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_7_sram;
wire [0:4] mux_tree_tapbuf_size17_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_8_sram;
wire [0:4] mux_tree_tapbuf_size17_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size17_9_sram;
wire [0:4] mux_tree_tapbuf_size17_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size17_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size17_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size23_0_sram;
wire [0:4] mux_tree_tapbuf_size23_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size23_1_sram;
wire [0:4] mux_tree_tapbuf_size23_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size23_2_sram;
wire [0:4] mux_tree_tapbuf_size23_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size23_3_sram;
wire [0:4] mux_tree_tapbuf_size23_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size23_4_sram;
wire [0:4] mux_tree_tapbuf_size23_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size23_5_sram;
wire [0:4] mux_tree_tapbuf_size23_5_sram_inv;
wire [0:0] mux_tree_tapbuf_size23_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size23_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size23_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size23_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size23_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size23_mem_5_ccff_tail;
wire [0:4] mux_tree_tapbuf_size24_0_sram;
wire [0:4] mux_tree_tapbuf_size24_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_10_sram;
wire [0:4] mux_tree_tapbuf_size24_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_11_sram;
wire [0:4] mux_tree_tapbuf_size24_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_12_sram;
wire [0:4] mux_tree_tapbuf_size24_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_13_sram;
wire [0:4] mux_tree_tapbuf_size24_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_14_sram;
wire [0:4] mux_tree_tapbuf_size24_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_15_sram;
wire [0:4] mux_tree_tapbuf_size24_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_16_sram;
wire [0:4] mux_tree_tapbuf_size24_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_17_sram;
wire [0:4] mux_tree_tapbuf_size24_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_18_sram;
wire [0:4] mux_tree_tapbuf_size24_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_19_sram;
wire [0:4] mux_tree_tapbuf_size24_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_1_sram;
wire [0:4] mux_tree_tapbuf_size24_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_20_sram;
wire [0:4] mux_tree_tapbuf_size24_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_21_sram;
wire [0:4] mux_tree_tapbuf_size24_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_22_sram;
wire [0:4] mux_tree_tapbuf_size24_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_23_sram;
wire [0:4] mux_tree_tapbuf_size24_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_24_sram;
wire [0:4] mux_tree_tapbuf_size24_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_25_sram;
wire [0:4] mux_tree_tapbuf_size24_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_26_sram;
wire [0:4] mux_tree_tapbuf_size24_26_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_27_sram;
wire [0:4] mux_tree_tapbuf_size24_27_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_28_sram;
wire [0:4] mux_tree_tapbuf_size24_28_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_29_sram;
wire [0:4] mux_tree_tapbuf_size24_29_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_2_sram;
wire [0:4] mux_tree_tapbuf_size24_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_30_sram;
wire [0:4] mux_tree_tapbuf_size24_30_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_31_sram;
wire [0:4] mux_tree_tapbuf_size24_31_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_32_sram;
wire [0:4] mux_tree_tapbuf_size24_32_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_33_sram;
wire [0:4] mux_tree_tapbuf_size24_33_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_34_sram;
wire [0:4] mux_tree_tapbuf_size24_34_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_35_sram;
wire [0:4] mux_tree_tapbuf_size24_35_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_36_sram;
wire [0:4] mux_tree_tapbuf_size24_36_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_37_sram;
wire [0:4] mux_tree_tapbuf_size24_37_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_38_sram;
wire [0:4] mux_tree_tapbuf_size24_38_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_39_sram;
wire [0:4] mux_tree_tapbuf_size24_39_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_3_sram;
wire [0:4] mux_tree_tapbuf_size24_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_40_sram;
wire [0:4] mux_tree_tapbuf_size24_40_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_41_sram;
wire [0:4] mux_tree_tapbuf_size24_41_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_42_sram;
wire [0:4] mux_tree_tapbuf_size24_42_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_43_sram;
wire [0:4] mux_tree_tapbuf_size24_43_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_44_sram;
wire [0:4] mux_tree_tapbuf_size24_44_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_45_sram;
wire [0:4] mux_tree_tapbuf_size24_45_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_46_sram;
wire [0:4] mux_tree_tapbuf_size24_46_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_47_sram;
wire [0:4] mux_tree_tapbuf_size24_47_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_48_sram;
wire [0:4] mux_tree_tapbuf_size24_48_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_49_sram;
wire [0:4] mux_tree_tapbuf_size24_49_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_4_sram;
wire [0:4] mux_tree_tapbuf_size24_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_50_sram;
wire [0:4] mux_tree_tapbuf_size24_50_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_51_sram;
wire [0:4] mux_tree_tapbuf_size24_51_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_52_sram;
wire [0:4] mux_tree_tapbuf_size24_52_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_53_sram;
wire [0:4] mux_tree_tapbuf_size24_53_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_54_sram;
wire [0:4] mux_tree_tapbuf_size24_54_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_55_sram;
wire [0:4] mux_tree_tapbuf_size24_55_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_56_sram;
wire [0:4] mux_tree_tapbuf_size24_56_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_57_sram;
wire [0:4] mux_tree_tapbuf_size24_57_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_58_sram;
wire [0:4] mux_tree_tapbuf_size24_58_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_59_sram;
wire [0:4] mux_tree_tapbuf_size24_59_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_5_sram;
wire [0:4] mux_tree_tapbuf_size24_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_60_sram;
wire [0:4] mux_tree_tapbuf_size24_60_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_61_sram;
wire [0:4] mux_tree_tapbuf_size24_61_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_62_sram;
wire [0:4] mux_tree_tapbuf_size24_62_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_63_sram;
wire [0:4] mux_tree_tapbuf_size24_63_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_64_sram;
wire [0:4] mux_tree_tapbuf_size24_64_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_65_sram;
wire [0:4] mux_tree_tapbuf_size24_65_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_6_sram;
wire [0:4] mux_tree_tapbuf_size24_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_7_sram;
wire [0:4] mux_tree_tapbuf_size24_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_8_sram;
wire [0:4] mux_tree_tapbuf_size24_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size24_9_sram;
wire [0:4] mux_tree_tapbuf_size24_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size24_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size24_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_4_sram;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_5_sram;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_6_sram;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_7_sram;
wire [0:2] mux_tree_tapbuf_size7_7_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail;
wire [0:3] mux_tree_tapbuf_size8_0_sram;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_100_sram;
wire [0:3] mux_tree_tapbuf_size8_100_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_101_sram;
wire [0:3] mux_tree_tapbuf_size8_101_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_102_sram;
wire [0:3] mux_tree_tapbuf_size8_102_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_103_sram;
wire [0:3] mux_tree_tapbuf_size8_103_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_104_sram;
wire [0:3] mux_tree_tapbuf_size8_104_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_105_sram;
wire [0:3] mux_tree_tapbuf_size8_105_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_106_sram;
wire [0:3] mux_tree_tapbuf_size8_106_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_107_sram;
wire [0:3] mux_tree_tapbuf_size8_107_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_10_sram;
wire [0:3] mux_tree_tapbuf_size8_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_11_sram;
wire [0:3] mux_tree_tapbuf_size8_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_12_sram;
wire [0:3] mux_tree_tapbuf_size8_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_13_sram;
wire [0:3] mux_tree_tapbuf_size8_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_14_sram;
wire [0:3] mux_tree_tapbuf_size8_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_15_sram;
wire [0:3] mux_tree_tapbuf_size8_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_16_sram;
wire [0:3] mux_tree_tapbuf_size8_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_17_sram;
wire [0:3] mux_tree_tapbuf_size8_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_18_sram;
wire [0:3] mux_tree_tapbuf_size8_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_19_sram;
wire [0:3] mux_tree_tapbuf_size8_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_1_sram;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_20_sram;
wire [0:3] mux_tree_tapbuf_size8_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_21_sram;
wire [0:3] mux_tree_tapbuf_size8_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_22_sram;
wire [0:3] mux_tree_tapbuf_size8_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_23_sram;
wire [0:3] mux_tree_tapbuf_size8_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_24_sram;
wire [0:3] mux_tree_tapbuf_size8_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_25_sram;
wire [0:3] mux_tree_tapbuf_size8_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_26_sram;
wire [0:3] mux_tree_tapbuf_size8_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_27_sram;
wire [0:3] mux_tree_tapbuf_size8_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_28_sram;
wire [0:3] mux_tree_tapbuf_size8_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_29_sram;
wire [0:3] mux_tree_tapbuf_size8_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_2_sram;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_30_sram;
wire [0:3] mux_tree_tapbuf_size8_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_31_sram;
wire [0:3] mux_tree_tapbuf_size8_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_32_sram;
wire [0:3] mux_tree_tapbuf_size8_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_33_sram;
wire [0:3] mux_tree_tapbuf_size8_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_34_sram;
wire [0:3] mux_tree_tapbuf_size8_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_35_sram;
wire [0:3] mux_tree_tapbuf_size8_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_36_sram;
wire [0:3] mux_tree_tapbuf_size8_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_37_sram;
wire [0:3] mux_tree_tapbuf_size8_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_38_sram;
wire [0:3] mux_tree_tapbuf_size8_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_39_sram;
wire [0:3] mux_tree_tapbuf_size8_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_3_sram;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_40_sram;
wire [0:3] mux_tree_tapbuf_size8_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_41_sram;
wire [0:3] mux_tree_tapbuf_size8_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_42_sram;
wire [0:3] mux_tree_tapbuf_size8_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_43_sram;
wire [0:3] mux_tree_tapbuf_size8_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_44_sram;
wire [0:3] mux_tree_tapbuf_size8_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_45_sram;
wire [0:3] mux_tree_tapbuf_size8_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_46_sram;
wire [0:3] mux_tree_tapbuf_size8_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_47_sram;
wire [0:3] mux_tree_tapbuf_size8_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_48_sram;
wire [0:3] mux_tree_tapbuf_size8_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_49_sram;
wire [0:3] mux_tree_tapbuf_size8_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_4_sram;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_50_sram;
wire [0:3] mux_tree_tapbuf_size8_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_51_sram;
wire [0:3] mux_tree_tapbuf_size8_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_52_sram;
wire [0:3] mux_tree_tapbuf_size8_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_53_sram;
wire [0:3] mux_tree_tapbuf_size8_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_54_sram;
wire [0:3] mux_tree_tapbuf_size8_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_55_sram;
wire [0:3] mux_tree_tapbuf_size8_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_56_sram;
wire [0:3] mux_tree_tapbuf_size8_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_57_sram;
wire [0:3] mux_tree_tapbuf_size8_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_58_sram;
wire [0:3] mux_tree_tapbuf_size8_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_59_sram;
wire [0:3] mux_tree_tapbuf_size8_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_5_sram;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_60_sram;
wire [0:3] mux_tree_tapbuf_size8_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_61_sram;
wire [0:3] mux_tree_tapbuf_size8_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_62_sram;
wire [0:3] mux_tree_tapbuf_size8_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_63_sram;
wire [0:3] mux_tree_tapbuf_size8_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_64_sram;
wire [0:3] mux_tree_tapbuf_size8_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_65_sram;
wire [0:3] mux_tree_tapbuf_size8_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_66_sram;
wire [0:3] mux_tree_tapbuf_size8_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_67_sram;
wire [0:3] mux_tree_tapbuf_size8_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_68_sram;
wire [0:3] mux_tree_tapbuf_size8_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_69_sram;
wire [0:3] mux_tree_tapbuf_size8_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_6_sram;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_70_sram;
wire [0:3] mux_tree_tapbuf_size8_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_71_sram;
wire [0:3] mux_tree_tapbuf_size8_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_72_sram;
wire [0:3] mux_tree_tapbuf_size8_72_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_73_sram;
wire [0:3] mux_tree_tapbuf_size8_73_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_74_sram;
wire [0:3] mux_tree_tapbuf_size8_74_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_75_sram;
wire [0:3] mux_tree_tapbuf_size8_75_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_76_sram;
wire [0:3] mux_tree_tapbuf_size8_76_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_77_sram;
wire [0:3] mux_tree_tapbuf_size8_77_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_78_sram;
wire [0:3] mux_tree_tapbuf_size8_78_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_79_sram;
wire [0:3] mux_tree_tapbuf_size8_79_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_7_sram;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_80_sram;
wire [0:3] mux_tree_tapbuf_size8_80_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_81_sram;
wire [0:3] mux_tree_tapbuf_size8_81_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_82_sram;
wire [0:3] mux_tree_tapbuf_size8_82_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_83_sram;
wire [0:3] mux_tree_tapbuf_size8_83_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_84_sram;
wire [0:3] mux_tree_tapbuf_size8_84_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_85_sram;
wire [0:3] mux_tree_tapbuf_size8_85_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_86_sram;
wire [0:3] mux_tree_tapbuf_size8_86_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_87_sram;
wire [0:3] mux_tree_tapbuf_size8_87_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_88_sram;
wire [0:3] mux_tree_tapbuf_size8_88_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_89_sram;
wire [0:3] mux_tree_tapbuf_size8_89_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_8_sram;
wire [0:3] mux_tree_tapbuf_size8_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_90_sram;
wire [0:3] mux_tree_tapbuf_size8_90_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_91_sram;
wire [0:3] mux_tree_tapbuf_size8_91_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_92_sram;
wire [0:3] mux_tree_tapbuf_size8_92_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_93_sram;
wire [0:3] mux_tree_tapbuf_size8_93_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_94_sram;
wire [0:3] mux_tree_tapbuf_size8_94_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_95_sram;
wire [0:3] mux_tree_tapbuf_size8_95_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_96_sram;
wire [0:3] mux_tree_tapbuf_size8_96_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_97_sram;
wire [0:3] mux_tree_tapbuf_size8_97_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_98_sram;
wire [0:3] mux_tree_tapbuf_size8_98_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_99_sram;
wire [0:3] mux_tree_tapbuf_size8_99_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_9_sram;
wire [0:3] mux_tree_tapbuf_size8_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_10_sram;
wire [0:3] mux_tree_tapbuf_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_11_sram;
wire [0:3] mux_tree_tapbuf_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_12_sram;
wire [0:3] mux_tree_tapbuf_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_13_sram;
wire [0:3] mux_tree_tapbuf_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_14_sram;
wire [0:3] mux_tree_tapbuf_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_15_sram;
wire [0:3] mux_tree_tapbuf_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_16_sram;
wire [0:3] mux_tree_tapbuf_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_17_sram;
wire [0:3] mux_tree_tapbuf_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_18_sram;
wire [0:3] mux_tree_tapbuf_size9_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_19_sram;
wire [0:3] mux_tree_tapbuf_size9_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_1_sram;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_20_sram;
wire [0:3] mux_tree_tapbuf_size9_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_21_sram;
wire [0:3] mux_tree_tapbuf_size9_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_22_sram;
wire [0:3] mux_tree_tapbuf_size9_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_23_sram;
wire [0:3] mux_tree_tapbuf_size9_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_24_sram;
wire [0:3] mux_tree_tapbuf_size9_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_25_sram;
wire [0:3] mux_tree_tapbuf_size9_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_26_sram;
wire [0:3] mux_tree_tapbuf_size9_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_27_sram;
wire [0:3] mux_tree_tapbuf_size9_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_2_sram;
wire [0:3] mux_tree_tapbuf_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_3_sram;
wire [0:3] mux_tree_tapbuf_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_4_sram;
wire [0:3] mux_tree_tapbuf_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_5_sram;
wire [0:3] mux_tree_tapbuf_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_6_sram;
wire [0:3] mux_tree_tapbuf_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_7_sram;
wire [0:3] mux_tree_tapbuf_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_8_sram;
wire [0:3] mux_tree_tapbuf_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_9_sram;
wire [0:3] mux_tree_tapbuf_size9_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[189] = chany_top_in[188];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[190] = chany_top_in[189];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[191] = chany_top_in[190];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[193] = chany_top_in[192];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[194] = chany_top_in[193];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[195] = chany_top_in[194];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[197] = chany_top_in[196];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[198] = chany_top_in[197];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[199] = chany_top_in[198];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[201] = chany_top_in[200];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[202] = chany_top_in[201];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[203] = chany_top_in[202];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[205] = chany_top_in[204];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[206] = chany_top_in[205];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[207] = chany_top_in[206];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[209] = chany_top_in[208];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[210] = chany_top_in[209];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[211] = chany_top_in[210];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[213] = chany_top_in[212];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[214] = chany_top_in[213];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[215] = chany_top_in[214];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[217] = chany_top_in[216];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[218] = chany_top_in[217];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[219] = chany_top_in[218];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[221] = chany_top_in[220];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[222] = chany_top_in[221];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[223] = chany_top_in[222];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[225] = chany_top_in[224];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[226] = chany_top_in[225];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[227] = chany_top_in[226];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[229] = chany_top_in[228];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[230] = chany_top_in[229];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[231] = chany_top_in[230];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[233] = chany_top_in[232];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[234] = chany_top_in[233];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[235] = chany_top_in[234];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[237] = chany_top_in[236];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[238] = chany_top_in[237];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[239] = chany_top_in[238];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[241] = chany_top_in[240];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[242] = chany_top_in[241];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[243] = chany_top_in[242];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[245] = chany_top_in[244];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[246] = chany_top_in[245];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[247] = chany_top_in[246];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[249] = chany_top_in[248];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[250] = chany_top_in[249];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[251] = chany_top_in[250];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[253] = chany_top_in[252];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[254] = chany_top_in[253];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[255] = chany_top_in[254];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[257] = chany_top_in[256];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[258] = chany_top_in[257];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[259] = chany_top_in[258];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[261] = chany_top_in[260];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[262] = chany_top_in[261];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[263] = chany_top_in[262];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[265] = chany_top_in[264];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[266] = chany_top_in[265];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[267] = chany_top_in[266];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[269] = chany_top_in[268];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[270] = chany_top_in[269];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[271] = chany_top_in[270];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[273] = chany_top_in[272];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[274] = chany_top_in[273];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[275] = chany_top_in[274];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[277] = chany_top_in[276];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[278] = chany_top_in[277];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[279] = chany_top_in[278];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[281] = chany_top_in[280];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[282] = chany_top_in[281];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[283] = chany_top_in[282];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 533 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 537 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 541 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 543 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 545 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 547 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 549 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 551 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 553 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 555 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 557 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 559 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 561 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 563 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 565 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 567 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 569 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 570 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 571 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 573 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 574 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 575 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 577 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 578 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 579 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 581 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 582 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 583 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 585 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 586 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 587 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 589 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 590 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 591 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 593 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 594 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 595 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 597 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 598 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 599 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 601 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 602 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 603 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 605 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[177] = chanx_right_in[176];
// ----- Local connection due to Wire 606 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[178] = chanx_right_in[177];
// ----- Local connection due to Wire 607 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[179] = chanx_right_in[178];
// ----- Local connection due to Wire 609 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[181] = chanx_right_in[180];
// ----- Local connection due to Wire 610 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[182] = chanx_right_in[181];
// ----- Local connection due to Wire 611 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[183] = chanx_right_in[182];
// ----- Local connection due to Wire 613 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[185] = chanx_right_in[184];
// ----- Local connection due to Wire 614 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[186] = chanx_right_in[185];
// ----- Local connection due to Wire 615 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[187] = chanx_right_in[186];
// ----- Local connection due to Wire 617 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[189] = chanx_right_in[188];
// ----- Local connection due to Wire 618 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[190] = chanx_right_in[189];
// ----- Local connection due to Wire 619 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[191] = chanx_right_in[190];
// ----- Local connection due to Wire 621 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[193] = chanx_right_in[192];
// ----- Local connection due to Wire 622 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[194] = chanx_right_in[193];
// ----- Local connection due to Wire 623 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[195] = chanx_right_in[194];
// ----- Local connection due to Wire 625 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[197] = chanx_right_in[196];
// ----- Local connection due to Wire 626 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[198] = chanx_right_in[197];
// ----- Local connection due to Wire 627 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[199] = chanx_right_in[198];
// ----- Local connection due to Wire 629 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[201] = chanx_right_in[200];
// ----- Local connection due to Wire 630 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[202] = chanx_right_in[201];
// ----- Local connection due to Wire 631 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[203] = chanx_right_in[202];
// ----- Local connection due to Wire 633 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[205] = chanx_right_in[204];
// ----- Local connection due to Wire 634 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[206] = chanx_right_in[205];
// ----- Local connection due to Wire 635 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[207] = chanx_right_in[206];
// ----- Local connection due to Wire 637 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[209] = chanx_right_in[208];
// ----- Local connection due to Wire 638 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[210] = chanx_right_in[209];
// ----- Local connection due to Wire 639 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[211] = chanx_right_in[210];
// ----- Local connection due to Wire 641 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[213] = chanx_right_in[212];
// ----- Local connection due to Wire 642 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[214] = chanx_right_in[213];
// ----- Local connection due to Wire 643 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[215] = chanx_right_in[214];
// ----- Local connection due to Wire 645 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[217] = chanx_right_in[216];
// ----- Local connection due to Wire 646 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[218] = chanx_right_in[217];
// ----- Local connection due to Wire 647 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[219] = chanx_right_in[218];
// ----- Local connection due to Wire 649 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[221] = chanx_right_in[220];
// ----- Local connection due to Wire 650 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[222] = chanx_right_in[221];
// ----- Local connection due to Wire 651 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[223] = chanx_right_in[222];
// ----- Local connection due to Wire 653 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[225] = chanx_right_in[224];
// ----- Local connection due to Wire 654 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[226] = chanx_right_in[225];
// ----- Local connection due to Wire 655 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[227] = chanx_right_in[226];
// ----- Local connection due to Wire 657 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[229] = chanx_right_in[228];
// ----- Local connection due to Wire 658 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[230] = chanx_right_in[229];
// ----- Local connection due to Wire 659 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[231] = chanx_right_in[230];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[233] = chanx_right_in[232];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[234] = chanx_right_in[233];
// ----- Local connection due to Wire 663 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[235] = chanx_right_in[234];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[237] = chanx_right_in[236];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[238] = chanx_right_in[237];
// ----- Local connection due to Wire 667 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[239] = chanx_right_in[238];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[241] = chanx_right_in[240];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[242] = chanx_right_in[241];
// ----- Local connection due to Wire 671 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[243] = chanx_right_in[242];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[245] = chanx_right_in[244];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[246] = chanx_right_in[245];
// ----- Local connection due to Wire 675 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[247] = chanx_right_in[246];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[249] = chanx_right_in[248];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[250] = chanx_right_in[249];
// ----- Local connection due to Wire 679 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[251] = chanx_right_in[250];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[253] = chanx_right_in[252];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[254] = chanx_right_in[253];
// ----- Local connection due to Wire 683 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[255] = chanx_right_in[254];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[257] = chanx_right_in[256];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[258] = chanx_right_in[257];
// ----- Local connection due to Wire 687 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[259] = chanx_right_in[258];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[261] = chanx_right_in[260];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[262] = chanx_right_in[261];
// ----- Local connection due to Wire 691 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[263] = chanx_right_in[262];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[265] = chanx_right_in[264];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[266] = chanx_right_in[265];
// ----- Local connection due to Wire 695 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[267] = chanx_right_in[266];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[269] = chanx_right_in[268];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[270] = chanx_right_in[269];
// ----- Local connection due to Wire 699 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[271] = chanx_right_in[270];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[273] = chanx_right_in[272];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[274] = chanx_right_in[273];
// ----- Local connection due to Wire 703 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[275] = chanx_right_in[274];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[277] = chanx_right_in[276];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[278] = chanx_right_in[277];
// ----- Local connection due to Wire 707 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[279] = chanx_right_in[278];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[281] = chanx_right_in[280];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[282] = chanx_right_in[281];
// ----- Local connection due to Wire 711 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[283] = chanx_right_in[282];
// ----- Local connection due to Wire 789 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 791 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 793 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 795 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 797 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 799 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 801 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 803 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 805 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 807 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 809 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 811 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 813 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 815 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 817 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 819 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 821 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 822 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 823 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 825 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 826 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 827 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 829 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 830 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 831 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 833 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 834 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 835 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 837 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 838 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 839 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 841 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 842 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 843 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 845 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 846 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 847 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 849 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 850 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 851 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 853 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 854 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 855 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 857 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 858 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 859 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 861 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 862 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 863 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 865 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 866 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 867 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 869 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 870 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 871 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 873 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 874 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 875 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 877 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 878 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 879 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 881 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 882 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 883 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 885 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 886 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 887 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 889 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 890 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 891 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 893 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 894 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 895 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 897 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 898 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 899 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 901 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 902 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 903 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 905 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 906 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 907 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 909 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 910 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 911 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 913 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 914 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 915 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 917 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 918 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 919 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 921 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 922 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 923 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 925 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 926 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 927 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 929 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 930 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 931 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 933 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 934 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 935 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 937 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 938 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 939 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 941 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 942 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 943 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 945 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 946 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 947 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 949 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 950 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 951 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 953 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 954 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 955 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 957 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 958 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 959 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 961 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 962 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 963 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 965 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 966 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 967 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 969 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 970 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 971 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 973 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 974 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 975 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 977 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[189] = chany_bottom_in[188];
// ----- Local connection due to Wire 978 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[190] = chany_bottom_in[189];
// ----- Local connection due to Wire 979 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[191] = chany_bottom_in[190];
// ----- Local connection due to Wire 981 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[193] = chany_bottom_in[192];
// ----- Local connection due to Wire 982 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[194] = chany_bottom_in[193];
// ----- Local connection due to Wire 983 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[195] = chany_bottom_in[194];
// ----- Local connection due to Wire 985 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[197] = chany_bottom_in[196];
// ----- Local connection due to Wire 986 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[198] = chany_bottom_in[197];
// ----- Local connection due to Wire 987 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[199] = chany_bottom_in[198];
// ----- Local connection due to Wire 989 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[201] = chany_bottom_in[200];
// ----- Local connection due to Wire 990 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[202] = chany_bottom_in[201];
// ----- Local connection due to Wire 991 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[203] = chany_bottom_in[202];
// ----- Local connection due to Wire 993 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[205] = chany_bottom_in[204];
// ----- Local connection due to Wire 994 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[206] = chany_bottom_in[205];
// ----- Local connection due to Wire 995 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[207] = chany_bottom_in[206];
// ----- Local connection due to Wire 997 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[209] = chany_bottom_in[208];
// ----- Local connection due to Wire 998 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[210] = chany_bottom_in[209];
// ----- Local connection due to Wire 999 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[211] = chany_bottom_in[210];
// ----- Local connection due to Wire 1001 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[213] = chany_bottom_in[212];
// ----- Local connection due to Wire 1002 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[214] = chany_bottom_in[213];
// ----- Local connection due to Wire 1003 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[215] = chany_bottom_in[214];
// ----- Local connection due to Wire 1005 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[217] = chany_bottom_in[216];
// ----- Local connection due to Wire 1006 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[218] = chany_bottom_in[217];
// ----- Local connection due to Wire 1007 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[219] = chany_bottom_in[218];
// ----- Local connection due to Wire 1009 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[221] = chany_bottom_in[220];
// ----- Local connection due to Wire 1010 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[222] = chany_bottom_in[221];
// ----- Local connection due to Wire 1011 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[223] = chany_bottom_in[222];
// ----- Local connection due to Wire 1013 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[225] = chany_bottom_in[224];
// ----- Local connection due to Wire 1014 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[226] = chany_bottom_in[225];
// ----- Local connection due to Wire 1015 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[227] = chany_bottom_in[226];
// ----- Local connection due to Wire 1017 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[229] = chany_bottom_in[228];
// ----- Local connection due to Wire 1018 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[230] = chany_bottom_in[229];
// ----- Local connection due to Wire 1019 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[231] = chany_bottom_in[230];
// ----- Local connection due to Wire 1021 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[233] = chany_bottom_in[232];
// ----- Local connection due to Wire 1022 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[234] = chany_bottom_in[233];
// ----- Local connection due to Wire 1023 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[235] = chany_bottom_in[234];
// ----- Local connection due to Wire 1025 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[237] = chany_bottom_in[236];
// ----- Local connection due to Wire 1026 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[238] = chany_bottom_in[237];
// ----- Local connection due to Wire 1027 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[239] = chany_bottom_in[238];
// ----- Local connection due to Wire 1029 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[241] = chany_bottom_in[240];
// ----- Local connection due to Wire 1030 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[242] = chany_bottom_in[241];
// ----- Local connection due to Wire 1031 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[243] = chany_bottom_in[242];
// ----- Local connection due to Wire 1033 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[245] = chany_bottom_in[244];
// ----- Local connection due to Wire 1034 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[246] = chany_bottom_in[245];
// ----- Local connection due to Wire 1035 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[247] = chany_bottom_in[246];
// ----- Local connection due to Wire 1037 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[249] = chany_bottom_in[248];
// ----- Local connection due to Wire 1038 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[250] = chany_bottom_in[249];
// ----- Local connection due to Wire 1039 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[251] = chany_bottom_in[250];
// ----- Local connection due to Wire 1041 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[253] = chany_bottom_in[252];
// ----- Local connection due to Wire 1042 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[254] = chany_bottom_in[253];
// ----- Local connection due to Wire 1043 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[255] = chany_bottom_in[254];
// ----- Local connection due to Wire 1045 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[257] = chany_bottom_in[256];
// ----- Local connection due to Wire 1046 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[258] = chany_bottom_in[257];
// ----- Local connection due to Wire 1047 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[259] = chany_bottom_in[258];
// ----- Local connection due to Wire 1049 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[261] = chany_bottom_in[260];
// ----- Local connection due to Wire 1050 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[262] = chany_bottom_in[261];
// ----- Local connection due to Wire 1051 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[263] = chany_bottom_in[262];
// ----- Local connection due to Wire 1053 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[265] = chany_bottom_in[264];
// ----- Local connection due to Wire 1054 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[266] = chany_bottom_in[265];
// ----- Local connection due to Wire 1055 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[267] = chany_bottom_in[266];
// ----- Local connection due to Wire 1057 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[269] = chany_bottom_in[268];
// ----- Local connection due to Wire 1058 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[270] = chany_bottom_in[269];
// ----- Local connection due to Wire 1059 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[271] = chany_bottom_in[270];
// ----- Local connection due to Wire 1061 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[273] = chany_bottom_in[272];
// ----- Local connection due to Wire 1062 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[274] = chany_bottom_in[273];
// ----- Local connection due to Wire 1063 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[275] = chany_bottom_in[274];
// ----- Local connection due to Wire 1065 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[277] = chany_bottom_in[276];
// ----- Local connection due to Wire 1066 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[278] = chany_bottom_in[277];
// ----- Local connection due to Wire 1067 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[279] = chany_bottom_in[278];
// ----- Local connection due to Wire 1069 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[281] = chany_bottom_in[280];
// ----- Local connection due to Wire 1070 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[282] = chany_bottom_in[281];
// ----- Local connection due to Wire 1071 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[283] = chany_bottom_in[282];
// ----- Local connection due to Wire 1076 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 1077 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 1078 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 1080 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 1081 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 1082 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 1084 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 1085 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 1086 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 1088 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 1089 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 1090 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 1092 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 1093 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 1094 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 1096 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 1097 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 1098 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 1100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 1101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 1102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 1104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 1105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 1106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 1108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 1109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 1110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 1112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 1113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 1114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 1116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 1117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 1118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 1120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 1121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 1122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 1124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 1125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 1126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 1128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 1129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 1130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 1132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 1133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 1134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 1136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 1137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 1138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 1140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 1141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 1142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 1144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 1145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 1146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 1148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 1149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 1150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 1152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 1153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 1154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 1156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 1157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 1158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 1160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 1161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 1162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 1164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 1165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 1166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 1168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 1169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 1170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 1172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 1173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 1174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 1176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 1177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 1178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 1180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 1181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 1182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 1184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 1185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 1186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 1188 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 1189 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 1190 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 1192 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 1193 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 1194 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 1196 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 1197 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 1198 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 1200 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 1201 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 1202 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 1204 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 1205 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 1206 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 1208 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 1209 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 1210 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 1212 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 1213 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 1214 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 1216 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 1217 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 1218 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 1220 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 1221 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 1222 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 1224 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 1225 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 1226 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 1228 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 1229 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 1230 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 1232 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 1233 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 1234 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 1236 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 1237 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 1238 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 1240 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 1241 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 1242 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 1244 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 1245 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 1246 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 1248 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 1249 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 1250 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- Local connection due to Wire 1252 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[177] = chanx_left_in[176];
// ----- Local connection due to Wire 1253 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[178] = chanx_left_in[177];
// ----- Local connection due to Wire 1254 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[179] = chanx_left_in[178];
// ----- Local connection due to Wire 1256 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[181] = chanx_left_in[180];
// ----- Local connection due to Wire 1257 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[182] = chanx_left_in[181];
// ----- Local connection due to Wire 1258 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[183] = chanx_left_in[182];
// ----- Local connection due to Wire 1260 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[185] = chanx_left_in[184];
// ----- Local connection due to Wire 1261 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[186] = chanx_left_in[185];
// ----- Local connection due to Wire 1262 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[187] = chanx_left_in[186];
// ----- Local connection due to Wire 1264 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[189] = chanx_left_in[188];
// ----- Local connection due to Wire 1265 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[190] = chanx_left_in[189];
// ----- Local connection due to Wire 1266 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[191] = chanx_left_in[190];
// ----- Local connection due to Wire 1268 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[193] = chanx_left_in[192];
// ----- Local connection due to Wire 1269 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[194] = chanx_left_in[193];
// ----- Local connection due to Wire 1270 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[195] = chanx_left_in[194];
// ----- Local connection due to Wire 1272 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[197] = chanx_left_in[196];
// ----- Local connection due to Wire 1273 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[198] = chanx_left_in[197];
// ----- Local connection due to Wire 1274 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[199] = chanx_left_in[198];
// ----- Local connection due to Wire 1276 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[201] = chanx_left_in[200];
// ----- Local connection due to Wire 1277 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[202] = chanx_left_in[201];
// ----- Local connection due to Wire 1278 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[203] = chanx_left_in[202];
// ----- Local connection due to Wire 1280 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[205] = chanx_left_in[204];
// ----- Local connection due to Wire 1281 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[206] = chanx_left_in[205];
// ----- Local connection due to Wire 1282 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[207] = chanx_left_in[206];
// ----- Local connection due to Wire 1284 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[209] = chanx_left_in[208];
// ----- Local connection due to Wire 1285 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[210] = chanx_left_in[209];
// ----- Local connection due to Wire 1286 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[211] = chanx_left_in[210];
// ----- Local connection due to Wire 1288 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[213] = chanx_left_in[212];
// ----- Local connection due to Wire 1289 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[214] = chanx_left_in[213];
// ----- Local connection due to Wire 1290 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[215] = chanx_left_in[214];
// ----- Local connection due to Wire 1292 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[217] = chanx_left_in[216];
// ----- Local connection due to Wire 1293 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[218] = chanx_left_in[217];
// ----- Local connection due to Wire 1294 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[219] = chanx_left_in[218];
// ----- Local connection due to Wire 1296 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[221] = chanx_left_in[220];
// ----- Local connection due to Wire 1297 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[222] = chanx_left_in[221];
// ----- Local connection due to Wire 1298 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[223] = chanx_left_in[222];
// ----- Local connection due to Wire 1300 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[225] = chanx_left_in[224];
// ----- Local connection due to Wire 1301 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[226] = chanx_left_in[225];
// ----- Local connection due to Wire 1302 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[227] = chanx_left_in[226];
// ----- Local connection due to Wire 1304 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[229] = chanx_left_in[228];
// ----- Local connection due to Wire 1305 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[230] = chanx_left_in[229];
// ----- Local connection due to Wire 1306 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[231] = chanx_left_in[230];
// ----- Local connection due to Wire 1308 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[233] = chanx_left_in[232];
// ----- Local connection due to Wire 1309 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[234] = chanx_left_in[233];
// ----- Local connection due to Wire 1310 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[235] = chanx_left_in[234];
// ----- Local connection due to Wire 1312 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[237] = chanx_left_in[236];
// ----- Local connection due to Wire 1313 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[238] = chanx_left_in[237];
// ----- Local connection due to Wire 1314 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[239] = chanx_left_in[238];
// ----- Local connection due to Wire 1316 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[241] = chanx_left_in[240];
// ----- Local connection due to Wire 1317 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[242] = chanx_left_in[241];
// ----- Local connection due to Wire 1318 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[243] = chanx_left_in[242];
// ----- Local connection due to Wire 1320 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[245] = chanx_left_in[244];
// ----- Local connection due to Wire 1321 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[246] = chanx_left_in[245];
// ----- Local connection due to Wire 1322 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[247] = chanx_left_in[246];
// ----- Local connection due to Wire 1324 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[249] = chanx_left_in[248];
// ----- Local connection due to Wire 1325 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[250] = chanx_left_in[249];
// ----- Local connection due to Wire 1326 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[251] = chanx_left_in[250];
// ----- Local connection due to Wire 1328 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[253] = chanx_left_in[252];
// ----- Local connection due to Wire 1329 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[254] = chanx_left_in[253];
// ----- Local connection due to Wire 1330 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[255] = chanx_left_in[254];
// ----- Local connection due to Wire 1332 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[257] = chanx_left_in[256];
// ----- Local connection due to Wire 1333 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[258] = chanx_left_in[257];
// ----- Local connection due to Wire 1334 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[259] = chanx_left_in[258];
// ----- Local connection due to Wire 1336 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[261] = chanx_left_in[260];
// ----- Local connection due to Wire 1337 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[262] = chanx_left_in[261];
// ----- Local connection due to Wire 1338 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[263] = chanx_left_in[262];
// ----- Local connection due to Wire 1340 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[265] = chanx_left_in[264];
// ----- Local connection due to Wire 1341 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[266] = chanx_left_in[265];
// ----- Local connection due to Wire 1342 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[267] = chanx_left_in[266];
// ----- Local connection due to Wire 1344 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[269] = chanx_left_in[268];
// ----- Local connection due to Wire 1345 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[270] = chanx_left_in[269];
// ----- Local connection due to Wire 1346 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[271] = chanx_left_in[270];
// ----- Local connection due to Wire 1348 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[273] = chanx_left_in[272];
// ----- Local connection due to Wire 1349 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[274] = chanx_left_in[273];
// ----- Local connection due to Wire 1350 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[275] = chanx_left_in[274];
// ----- Local connection due to Wire 1352 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[277] = chanx_left_in[276];
// ----- Local connection due to Wire 1353 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[278] = chanx_left_in[277];
// ----- Local connection due to Wire 1354 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[279] = chanx_left_in[278];
// ----- Local connection due to Wire 1356 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[281] = chanx_left_in[280];
// ----- Local connection due to Wire 1357 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[282] = chanx_left_in[281];
// ----- Local connection due to Wire 1358 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[283] = chanx_left_in[282];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size24 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[97], chanx_right_in[193], chanx_left_in[0], chanx_left_in[3], chanx_left_in[96], chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size24_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_0_sram_inv[0:4]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size24 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[6], chanx_right_in[23], chanx_right_in[102], chanx_right_in[198], chanx_left_in[90], chanx_left_in[186], chanx_left_in[275], chanx_left_in[282]}),
		.sram(mux_tree_tapbuf_size24_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_1_sram_inv[0:4]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size24 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[104], chanx_right_in[200], chanx_left_in[89], chanx_left_in[185], chanx_left_in[271], chanx_left_in[281]}),
		.sram(mux_tree_tapbuf_size24_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_2_sram_inv[0:4]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size24 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[9], chanx_right_in[31], chanx_right_in[105], chanx_right_in[201], chanx_left_in[88], chanx_left_in[184], chanx_left_in[267], chanx_left_in[280]}),
		.sram(mux_tree_tapbuf_size24_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_3_sram_inv[0:4]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size24 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[10], chanx_right_in[35], chanx_right_in[106], chanx_right_in[202], chanx_left_in[86], chanx_left_in[182], chanx_left_in[263], chanx_left_in[278]}),
		.sram(mux_tree_tapbuf_size24_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_4_sram_inv[0:4]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size24 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[12], chanx_right_in[39], chanx_right_in[108], chanx_right_in[204], chanx_left_in[85], chanx_left_in[181], chanx_left_in[259], chanx_left_in[277]}),
		.sram(mux_tree_tapbuf_size24_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_5_sram_inv[0:4]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size24 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[13], chanx_right_in[43], chanx_right_in[109], chanx_right_in[205], chanx_left_in[84], chanx_left_in[180], chanx_left_in[255], chanx_left_in[276]}),
		.sram(mux_tree_tapbuf_size24_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_6_sram_inv[0:4]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size24 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[14], chanx_right_in[47], chanx_right_in[110], chanx_right_in[206], chanx_left_in[82], chanx_left_in[178], chanx_left_in[251], chanx_left_in[274]}),
		.sram(mux_tree_tapbuf_size24_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_7_sram_inv[0:4]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size24 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[16], chanx_right_in[51], chanx_right_in[112], chanx_right_in[208], chanx_left_in[81], chanx_left_in[177], chanx_left_in[247], chanx_left_in[273]}),
		.sram(mux_tree_tapbuf_size24_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_8_sram_inv[0:4]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size24 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[17], chanx_right_in[55], chanx_right_in[113], chanx_right_in[209], chanx_left_in[80], chanx_left_in[176], chanx_left_in[243], chanx_left_in[272]}),
		.sram(mux_tree_tapbuf_size24_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_9_sram_inv[0:4]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size24 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[18], chanx_right_in[59], chanx_right_in[114], chanx_right_in[210], chanx_left_in[78], chanx_left_in[174], chanx_left_in[239], chanx_left_in[270]}),
		.sram(mux_tree_tapbuf_size24_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_10_sram_inv[0:4]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size24 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[20], chanx_right_in[63], chanx_right_in[116], chanx_right_in[212], chanx_left_in[77], chanx_left_in[173], chanx_left_in[235], chanx_left_in[269]}),
		.sram(mux_tree_tapbuf_size24_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_11_sram_inv[0:4]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size24 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[21], chanx_right_in[67], chanx_right_in[117], chanx_right_in[213], chanx_left_in[76], chanx_left_in[172], chanx_left_in[231], chanx_left_in[268]}),
		.sram(mux_tree_tapbuf_size24_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_12_sram_inv[0:4]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size24 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[22], chanx_right_in[71], chanx_right_in[118], chanx_right_in[214], chanx_left_in[74], chanx_left_in[170], chanx_left_in[227], chanx_left_in[266]}),
		.sram(mux_tree_tapbuf_size24_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_13_sram_inv[0:4]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size24 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[24], chanx_right_in[75], chanx_right_in[120], chanx_right_in[216], chanx_left_in[73], chanx_left_in[169], chanx_left_in[223], chanx_left_in[265]}),
		.sram(mux_tree_tapbuf_size24_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_14_sram_inv[0:4]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size24 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[25], chanx_right_in[79], chanx_right_in[121], chanx_right_in[217], chanx_left_in[72], chanx_left_in[168], chanx_left_in[219], chanx_left_in[264]}),
		.sram(mux_tree_tapbuf_size24_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_15_sram_inv[0:4]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size24 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[26], chanx_right_in[83], chanx_right_in[122], chanx_right_in[218], chanx_left_in[70], chanx_left_in[166], chanx_left_in[215], chanx_left_in[262]}),
		.sram(mux_tree_tapbuf_size24_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_16_sram_inv[0:4]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size24 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[28], chanx_right_in[87], chanx_right_in[124], chanx_right_in[220], chanx_left_in[69], chanx_left_in[165], chanx_left_in[211], chanx_left_in[261]}),
		.sram(mux_tree_tapbuf_size24_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_17_sram_inv[0:4]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size24 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[29], chanx_right_in[91], chanx_right_in[125], chanx_right_in[221], chanx_left_in[68], chanx_left_in[164], chanx_left_in[207], chanx_left_in[260]}),
		.sram(mux_tree_tapbuf_size24_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_18_sram_inv[0:4]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size24 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[30], chanx_right_in[95], chanx_right_in[126], chanx_right_in[222], chanx_left_in[66], chanx_left_in[162], chanx_left_in[203], chanx_left_in[258]}),
		.sram(mux_tree_tapbuf_size24_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_19_sram_inv[0:4]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size24 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[32], chanx_right_in[99], chanx_right_in[128], chanx_right_in[224], chanx_left_in[65], chanx_left_in[161], chanx_left_in[199], chanx_left_in[257]}),
		.sram(mux_tree_tapbuf_size24_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_20_sram_inv[0:4]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size24 mux_top_track_192 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[33], chanx_right_in[103], chanx_right_in[129], chanx_right_in[225], chanx_left_in[64], chanx_left_in[160], chanx_left_in[195], chanx_left_in[256]}),
		.sram(mux_tree_tapbuf_size24_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_21_sram_inv[0:4]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size24 mux_top_track_200 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[34], chanx_right_in[107], chanx_right_in[130], chanx_right_in[226], chanx_left_in[62], chanx_left_in[158], chanx_left_in[191], chanx_left_in[254]}),
		.sram(mux_tree_tapbuf_size24_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_22_sram_inv[0:4]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size24 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[36], chanx_right_in[111], chanx_right_in[132], chanx_right_in[228], chanx_left_in[61], chanx_left_in[157], chanx_left_in[187], chanx_left_in[253]}),
		.sram(mux_tree_tapbuf_size24_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_23_sram_inv[0:4]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size24 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[37], chanx_right_in[115], chanx_right_in[133], chanx_right_in[229], chanx_left_in[60], chanx_left_in[156], chanx_left_in[183], chanx_left_in[252]}),
		.sram(mux_tree_tapbuf_size24_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_24_sram_inv[0:4]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size24 mux_top_track_224 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[38], chanx_right_in[119], chanx_right_in[134], chanx_right_in[230], chanx_left_in[58], chanx_left_in[154], chanx_left_in[179], chanx_left_in[250]}),
		.sram(mux_tree_tapbuf_size24_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_25_sram_inv[0:4]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size24 mux_top_track_232 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[40], chanx_right_in[123], chanx_right_in[136], chanx_right_in[232], chanx_left_in[57], chanx_left_in[153], chanx_left_in[175], chanx_left_in[249]}),
		.sram(mux_tree_tapbuf_size24_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_26_sram_inv[0:4]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size24 mux_top_track_240 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[41], chanx_right_in[127], chanx_right_in[137], chanx_right_in[233], chanx_left_in[56], chanx_left_in[152], chanx_left_in[171], chanx_left_in[248]}),
		.sram(mux_tree_tapbuf_size24_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_27_sram_inv[0:4]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size24 mux_top_track_248 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[42], chanx_right_in[131], chanx_right_in[138], chanx_right_in[234], chanx_left_in[54], chanx_left_in[150], chanx_left_in[167], chanx_left_in[246]}),
		.sram(mux_tree_tapbuf_size24_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_28_sram_inv[0:4]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size24 mux_top_track_256 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[44], chanx_right_in[135], chanx_right_in[140], chanx_right_in[236], chanx_left_in[53], chanx_left_in[149], chanx_left_in[163], chanx_left_in[245]}),
		.sram(mux_tree_tapbuf_size24_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_29_sram_inv[0:4]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size24 mux_top_track_264 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[45], chanx_right_in[139], chanx_right_in[141], chanx_right_in[237], chanx_left_in[52], chanx_left_in[148], chanx_left_in[159], chanx_left_in[244]}),
		.sram(mux_tree_tapbuf_size24_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_30_sram_inv[0:4]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size24 mux_top_track_272 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[46], chanx_right_in[142:143], chanx_right_in[238], chanx_left_in[50], chanx_left_in[146], chanx_left_in[155], chanx_left_in[242]}),
		.sram(mux_tree_tapbuf_size24_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_31_sram_inv[0:4]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size24 mux_top_track_280 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[48], chanx_right_in[144], chanx_right_in[147], chanx_right_in[240], chanx_left_in[49], chanx_left_in[145], chanx_left_in[151], chanx_left_in[241]}),
		.sram(mux_tree_tapbuf_size24_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_32_sram_inv[0:4]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size24 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[49], chanx_right_in[145], chanx_right_in[151], chanx_right_in[241], chanx_left_in[48], chanx_left_in[144], chanx_left_in[147], chanx_left_in[240]}),
		.sram(mux_tree_tapbuf_size24_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_33_sram_inv[0:4]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size24 mux_top_track_296 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[50], chanx_right_in[146], chanx_right_in[155], chanx_right_in[242], chanx_left_in[46], chanx_left_in[142:143], chanx_left_in[238]}),
		.sram(mux_tree_tapbuf_size24_34_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_34_sram_inv[0:4]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size24 mux_top_track_304 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[52], chanx_right_in[148], chanx_right_in[159], chanx_right_in[244], chanx_left_in[45], chanx_left_in[139], chanx_left_in[141], chanx_left_in[237]}),
		.sram(mux_tree_tapbuf_size24_35_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_35_sram_inv[0:4]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size24 mux_top_track_312 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[53], chanx_right_in[149], chanx_right_in[163], chanx_right_in[245], chanx_left_in[44], chanx_left_in[135], chanx_left_in[140], chanx_left_in[236]}),
		.sram(mux_tree_tapbuf_size24_36_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_36_sram_inv[0:4]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size24 mux_top_track_320 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[54], chanx_right_in[150], chanx_right_in[167], chanx_right_in[246], chanx_left_in[42], chanx_left_in[131], chanx_left_in[138], chanx_left_in[234]}),
		.sram(mux_tree_tapbuf_size24_37_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_37_sram_inv[0:4]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size24 mux_top_track_328 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[56], chanx_right_in[152], chanx_right_in[171], chanx_right_in[248], chanx_left_in[41], chanx_left_in[127], chanx_left_in[137], chanx_left_in[233]}),
		.sram(mux_tree_tapbuf_size24_38_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_38_sram_inv[0:4]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size24 mux_top_track_336 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[57], chanx_right_in[153], chanx_right_in[175], chanx_right_in[249], chanx_left_in[40], chanx_left_in[123], chanx_left_in[136], chanx_left_in[232]}),
		.sram(mux_tree_tapbuf_size24_39_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_39_sram_inv[0:4]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size24 mux_top_track_344 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[58], chanx_right_in[154], chanx_right_in[179], chanx_right_in[250], chanx_left_in[38], chanx_left_in[119], chanx_left_in[134], chanx_left_in[230]}),
		.sram(mux_tree_tapbuf_size24_40_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_40_sram_inv[0:4]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size24 mux_top_track_352 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[60], chanx_right_in[156], chanx_right_in[183], chanx_right_in[252], chanx_left_in[37], chanx_left_in[115], chanx_left_in[133], chanx_left_in[229]}),
		.sram(mux_tree_tapbuf_size24_41_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_41_sram_inv[0:4]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size24 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[61], chanx_right_in[157], chanx_right_in[187], chanx_right_in[253], chanx_left_in[36], chanx_left_in[111], chanx_left_in[132], chanx_left_in[228]}),
		.sram(mux_tree_tapbuf_size24_42_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_42_sram_inv[0:4]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size24 mux_top_track_368 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[62], chanx_right_in[158], chanx_right_in[191], chanx_right_in[254], chanx_left_in[34], chanx_left_in[107], chanx_left_in[130], chanx_left_in[226]}),
		.sram(mux_tree_tapbuf_size24_43_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_43_sram_inv[0:4]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size24 mux_top_track_376 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[64], chanx_right_in[160], chanx_right_in[195], chanx_right_in[256], chanx_left_in[33], chanx_left_in[103], chanx_left_in[129], chanx_left_in[225]}),
		.sram(mux_tree_tapbuf_size24_44_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_44_sram_inv[0:4]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size24 mux_top_track_384 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[65], chanx_right_in[161], chanx_right_in[199], chanx_right_in[257], chanx_left_in[32], chanx_left_in[99], chanx_left_in[128], chanx_left_in[224]}),
		.sram(mux_tree_tapbuf_size24_45_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_45_sram_inv[0:4]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size24 mux_top_track_392 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[66], chanx_right_in[162], chanx_right_in[203], chanx_right_in[258], chanx_left_in[30], chanx_left_in[95], chanx_left_in[126], chanx_left_in[222]}),
		.sram(mux_tree_tapbuf_size24_46_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_46_sram_inv[0:4]),
		.out(chany_top_out[196]));

	mux_tree_tapbuf_size24 mux_top_track_400 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[68], chanx_right_in[164], chanx_right_in[207], chanx_right_in[260], chanx_left_in[29], chanx_left_in[91], chanx_left_in[125], chanx_left_in[221]}),
		.sram(mux_tree_tapbuf_size24_47_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_47_sram_inv[0:4]),
		.out(chany_top_out[200]));

	mux_tree_tapbuf_size24 mux_top_track_408 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[69], chanx_right_in[165], chanx_right_in[211], chanx_right_in[261], chanx_left_in[28], chanx_left_in[87], chanx_left_in[124], chanx_left_in[220]}),
		.sram(mux_tree_tapbuf_size24_48_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_48_sram_inv[0:4]),
		.out(chany_top_out[204]));

	mux_tree_tapbuf_size24 mux_top_track_416 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[70], chanx_right_in[166], chanx_right_in[215], chanx_right_in[262], chanx_left_in[26], chanx_left_in[83], chanx_left_in[122], chanx_left_in[218]}),
		.sram(mux_tree_tapbuf_size24_49_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_49_sram_inv[0:4]),
		.out(chany_top_out[208]));

	mux_tree_tapbuf_size24 mux_top_track_424 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[72], chanx_right_in[168], chanx_right_in[219], chanx_right_in[264], chanx_left_in[25], chanx_left_in[79], chanx_left_in[121], chanx_left_in[217]}),
		.sram(mux_tree_tapbuf_size24_50_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_50_sram_inv[0:4]),
		.out(chany_top_out[212]));

	mux_tree_tapbuf_size24 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[73], chanx_right_in[169], chanx_right_in[223], chanx_right_in[265], chanx_left_in[24], chanx_left_in[75], chanx_left_in[120], chanx_left_in[216]}),
		.sram(mux_tree_tapbuf_size24_51_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_51_sram_inv[0:4]),
		.out(chany_top_out[216]));

	mux_tree_tapbuf_size24 mux_top_track_440 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[74], chanx_right_in[170], chanx_right_in[227], chanx_right_in[266], chanx_left_in[22], chanx_left_in[71], chanx_left_in[118], chanx_left_in[214]}),
		.sram(mux_tree_tapbuf_size24_52_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_52_sram_inv[0:4]),
		.out(chany_top_out[220]));

	mux_tree_tapbuf_size24 mux_top_track_448 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[76], chanx_right_in[172], chanx_right_in[231], chanx_right_in[268], chanx_left_in[21], chanx_left_in[67], chanx_left_in[117], chanx_left_in[213]}),
		.sram(mux_tree_tapbuf_size24_53_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_53_sram_inv[0:4]),
		.out(chany_top_out[224]));

	mux_tree_tapbuf_size24 mux_top_track_456 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[77], chanx_right_in[173], chanx_right_in[235], chanx_right_in[269], chanx_left_in[20], chanx_left_in[63], chanx_left_in[116], chanx_left_in[212]}),
		.sram(mux_tree_tapbuf_size24_54_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_54_sram_inv[0:4]),
		.out(chany_top_out[228]));

	mux_tree_tapbuf_size24 mux_top_track_464 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[78], chanx_right_in[174], chanx_right_in[239], chanx_right_in[270], chanx_left_in[18], chanx_left_in[59], chanx_left_in[114], chanx_left_in[210]}),
		.sram(mux_tree_tapbuf_size24_55_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_55_sram_inv[0:4]),
		.out(chany_top_out[232]));

	mux_tree_tapbuf_size24 mux_top_track_472 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[80], chanx_right_in[176], chanx_right_in[243], chanx_right_in[272], chanx_left_in[17], chanx_left_in[55], chanx_left_in[113], chanx_left_in[209]}),
		.sram(mux_tree_tapbuf_size24_56_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_56_sram_inv[0:4]),
		.out(chany_top_out[236]));

	mux_tree_tapbuf_size24 mux_top_track_480 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[81], chanx_right_in[177], chanx_right_in[247], chanx_right_in[273], chanx_left_in[16], chanx_left_in[51], chanx_left_in[112], chanx_left_in[208]}),
		.sram(mux_tree_tapbuf_size24_57_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_57_sram_inv[0:4]),
		.out(chany_top_out[240]));

	mux_tree_tapbuf_size24 mux_top_track_488 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[82], chanx_right_in[178], chanx_right_in[251], chanx_right_in[274], chanx_left_in[14], chanx_left_in[47], chanx_left_in[110], chanx_left_in[206]}),
		.sram(mux_tree_tapbuf_size24_58_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_58_sram_inv[0:4]),
		.out(chany_top_out[244]));

	mux_tree_tapbuf_size24 mux_top_track_496 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[84], chanx_right_in[180], chanx_right_in[255], chanx_right_in[276], chanx_left_in[13], chanx_left_in[43], chanx_left_in[109], chanx_left_in[205]}),
		.sram(mux_tree_tapbuf_size24_59_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_59_sram_inv[0:4]),
		.out(chany_top_out[248]));

	mux_tree_tapbuf_size24 mux_top_track_504 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_64_, chanx_right_in[85], chanx_right_in[181], chanx_right_in[259], chanx_right_in[277], chanx_left_in[12], chanx_left_in[39], chanx_left_in[108], chanx_left_in[204]}),
		.sram(mux_tree_tapbuf_size24_60_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_60_sram_inv[0:4]),
		.out(chany_top_out[252]));

	mux_tree_tapbuf_size24 mux_top_track_512 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[86], chanx_right_in[182], chanx_right_in[263], chanx_right_in[278], chanx_left_in[10], chanx_left_in[35], chanx_left_in[106], chanx_left_in[202]}),
		.sram(mux_tree_tapbuf_size24_61_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_61_sram_inv[0:4]),
		.out(chany_top_out[256]));

	mux_tree_tapbuf_size24 mux_top_track_520 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[88], chanx_right_in[184], chanx_right_in[267], chanx_right_in[280], chanx_left_in[9], chanx_left_in[31], chanx_left_in[105], chanx_left_in[201]}),
		.sram(mux_tree_tapbuf_size24_62_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_62_sram_inv[0:4]),
		.out(chany_top_out[260]));

	mux_tree_tapbuf_size24 mux_top_track_528 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[89], chanx_right_in[185], chanx_right_in[271], chanx_right_in[281], chanx_left_in[8], chanx_left_in[27], chanx_left_in[104], chanx_left_in[200]}),
		.sram(mux_tree_tapbuf_size24_63_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_63_sram_inv[0:4]),
		.out(chany_top_out[264]));

	mux_tree_tapbuf_size24 mux_top_track_536 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_66_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_68_, chanx_right_in[90], chanx_right_in[186], chanx_right_in[275], chanx_right_in[282], chanx_left_in[6], chanx_left_in[23], chanx_left_in[102], chanx_left_in[198]}),
		.sram(mux_tree_tapbuf_size24_64_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_64_sram_inv[0:4]),
		.out(chany_top_out[268]));

	mux_tree_tapbuf_size24 mux_top_track_568 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_2_, chanx_right_in[0], chanx_right_in[3], chanx_right_in[96], chanx_right_in[192], chanx_left_in[1], chanx_left_in[7], chanx_left_in[97], chanx_left_in[193]}),
		.sram(mux_tree_tapbuf_size24_65_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size24_65_sram_inv[0:4]),
		.out(chany_top_out[284]));

	mux_tree_tapbuf_size24_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size24_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_0_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_1_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_2_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_3_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_4_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_5_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_6_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_7_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_8_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_9_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_10_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_11_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_12_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_13_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_14_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_15_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_16_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_17_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_18_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_19_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_20_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_21_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_22_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_23_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_24_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_25_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_26_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_27_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_28_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_29_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_30_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_31_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_32_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_33_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_34_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_34_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_35_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_35_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_36_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_36_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_37_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_37_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_38_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_38_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_39_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_39_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_40_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_40_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_41_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_41_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_42_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_42_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_43_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_43_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_44_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_44_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_45_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_45_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_46_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_46_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_47_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_47_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_48_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_48_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_49_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_49_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_50_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_50_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_51_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_51_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_52_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_52_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_53_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_53_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_54_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_54_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_55_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_55_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_56_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_56_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_57_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_57_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_58_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_58_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_59_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_59_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_60_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_60_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_61_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_61_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_62_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_62_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_63_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_63_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_64_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_64_sram_inv[0:4]));

	mux_tree_tapbuf_size24_mem mem_top_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size24_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size24_65_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size24_65_sram_inv[0:4]));

	mux_tree_tapbuf_size23 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_36_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_54_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_63_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_65_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[98], chanx_right_in[194], chanx_left_in[94], chanx_left_in[190], chanx_left_in[284]}),
		.sram(mux_tree_tapbuf_size23_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_0_sram_inv[0:4]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size23 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_46_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_55_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_64_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_39_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_48_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_66_, chanx_right_in[4], chanx_right_in[15], chanx_right_in[100], chanx_right_in[196], chanx_left_in[93], chanx_left_in[189], chanx_left_in[283]}),
		.sram(mux_tree_tapbuf_size23_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_1_sram_inv[0:4]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size23 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_38_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_47_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_56_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_67_, chanx_right_in[5], chanx_right_in[19], chanx_right_in[101], chanx_right_in[197], chanx_left_in[92], chanx_left_in[188], chanx_left_in[279]}),
		.sram(mux_tree_tapbuf_size23_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_2_sram_inv[0:4]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size23 mux_top_track_544 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_40_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_58_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_67_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_69_, chanx_right_in[92], chanx_right_in[188], chanx_right_in[279], chanx_left_in[5], chanx_left_in[19], chanx_left_in[101], chanx_left_in[197]}),
		.sram(mux_tree_tapbuf_size23_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_3_sram_inv[0:4]),
		.out(chany_top_out[272]));

	mux_tree_tapbuf_size23 mux_top_track_552 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_50_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_59_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_68_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_43_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_52_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_0_, chanx_right_in[93], chanx_right_in[189], chanx_right_in[283], chanx_left_in[4], chanx_left_in[15], chanx_left_in[100], chanx_left_in[196]}),
		.sram(mux_tree_tapbuf_size23_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_4_sram_inv[0:4]),
		.out(chany_top_out[276]));

	mux_tree_tapbuf_size23 mux_top_track_560 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_42_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_51_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_60_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_3_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_35_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_44_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_4_62_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_1_, chanx_right_in[94], chanx_right_in[190], chanx_right_in[284], chanx_left_in[2], chanx_left_in[11], chanx_left_in[98], chanx_left_in[194]}),
		.sram(mux_tree_tapbuf_size23_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size23_5_sram_inv[0:4]),
		.out(chany_top_out[280]));

	mux_tree_tapbuf_size23_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_0_sram_inv[0:4]));

	mux_tree_tapbuf_size23_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_1_sram_inv[0:4]));

	mux_tree_tapbuf_size23_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_2_sram_inv[0:4]));

	mux_tree_tapbuf_size23_mem mem_top_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_3_sram_inv[0:4]));

	mux_tree_tapbuf_size23_mem mem_top_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_4_sram_inv[0:4]));

	mux_tree_tapbuf_size23_mem mem_top_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size23_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size23_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size23_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size23_5_sram_inv[0:4]));

	mux_tree_tapbuf_size15 mux_right_track_0 (
		.in({chany_top_in[94], chany_top_in[190], chany_top_in[284], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[93], chany_bottom_in[189], chany_bottom_in[283]}),
		.sram(mux_tree_tapbuf_size15_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size15 mux_right_track_560 (
		.in({chany_top_in[92], chany_top_in[188], chany_top_in[279], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[96], chany_bottom_in[192]}),
		.sram(mux_tree_tapbuf_size15_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_1_sram_inv[0:3]),
		.out(chanx_right_out[280]));

	mux_tree_tapbuf_size15_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size24_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_0_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_right_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_1_sram_inv[0:3]));

	mux_tree_tapbuf_size16 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[96], chany_top_in[192], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[92], chany_bottom_in[188], chany_bottom_in[279]}),
		.sram(mux_tree_tapbuf_size16_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_0_sram_inv[0:4]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size16 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[98], chany_top_in[194], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[89], chany_bottom_in[185], chany_bottom_in[271], chany_bottom_in[281]}),
		.sram(mux_tree_tapbuf_size16_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_1_sram_inv[0:4]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size16 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[100], chany_top_in[196], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[88], chany_bottom_in[184], chany_bottom_in[267], chany_bottom_in[280]}),
		.sram(mux_tree_tapbuf_size16_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_2_sram_inv[0:4]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size16 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[101], chany_top_in[197], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[86], chany_bottom_in[182], chany_bottom_in[263], chany_bottom_in[278]}),
		.sram(mux_tree_tapbuf_size16_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_3_sram_inv[0:4]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size16 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[102], chany_top_in[198], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[85], chany_bottom_in[181], chany_bottom_in[259], chany_bottom_in[277]}),
		.sram(mux_tree_tapbuf_size16_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_4_sram_inv[0:4]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size16 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[104], chany_top_in[200], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[84], chany_bottom_in[180], chany_bottom_in[255], chany_bottom_in[276]}),
		.sram(mux_tree_tapbuf_size16_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_5_sram_inv[0:4]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size16 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[105], chany_top_in[201], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[82], chany_bottom_in[178], chany_bottom_in[251], chany_bottom_in[274]}),
		.sram(mux_tree_tapbuf_size16_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_6_sram_inv[0:4]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size16 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[110], chany_top_in[206], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[77], chany_bottom_in[173], chany_bottom_in[235], chany_bottom_in[269]}),
		.sram(mux_tree_tapbuf_size16_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_7_sram_inv[0:4]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size16 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[112], chany_top_in[208], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[76], chany_bottom_in[172], chany_bottom_in[231], chany_bottom_in[268]}),
		.sram(mux_tree_tapbuf_size16_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_8_sram_inv[0:4]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size16 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[113], chany_top_in[209], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[74], chany_bottom_in[170], chany_bottom_in[227], chany_bottom_in[266]}),
		.sram(mux_tree_tapbuf_size16_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_9_sram_inv[0:4]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size16 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[114], chany_top_in[210], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[73], chany_bottom_in[169], chany_bottom_in[223], chany_bottom_in[265]}),
		.sram(mux_tree_tapbuf_size16_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_10_sram_inv[0:4]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size16 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[116], chany_top_in[212], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[72], chany_bottom_in[168], chany_bottom_in[219], chany_bottom_in[264]}),
		.sram(mux_tree_tapbuf_size16_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_11_sram_inv[0:4]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size16 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[117], chany_top_in[213], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[70], chany_bottom_in[166], chany_bottom_in[215], chany_bottom_in[262]}),
		.sram(mux_tree_tapbuf_size16_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_12_sram_inv[0:4]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size16 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[122], chany_top_in[218], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[65], chany_bottom_in[161], chany_bottom_in[199], chany_bottom_in[257]}),
		.sram(mux_tree_tapbuf_size16_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_13_sram_inv[0:4]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size16 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[124], chany_top_in[220], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[64], chany_bottom_in[160], chany_bottom_in[195], chany_bottom_in[256]}),
		.sram(mux_tree_tapbuf_size16_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_14_sram_inv[0:4]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size16 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[125], chany_top_in[221], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[62], chany_bottom_in[158], chany_bottom_in[191], chany_bottom_in[254]}),
		.sram(mux_tree_tapbuf_size16_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_15_sram_inv[0:4]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size16 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[95], chany_top_in[126], chany_top_in[222], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[61], chany_bottom_in[157], chany_bottom_in[187], chany_bottom_in[253]}),
		.sram(mux_tree_tapbuf_size16_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_16_sram_inv[0:4]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size16 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[99], chany_top_in[128], chany_top_in[224], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[60], chany_bottom_in[156], chany_bottom_in[183], chany_bottom_in[252]}),
		.sram(mux_tree_tapbuf_size16_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_17_sram_inv[0:4]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size16 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[103], chany_top_in[129], chany_top_in[225], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[58], chany_bottom_in[154], chany_bottom_in[179], chany_bottom_in[250]}),
		.sram(mux_tree_tapbuf_size16_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_18_sram_inv[0:4]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size16 mux_right_track_240 (
		.in({chany_top_in[38], chany_top_in[119], chany_top_in[134], chany_top_in[230], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[53], chany_bottom_in[149], chany_bottom_in[163], chany_bottom_in[245]}),
		.sram(mux_tree_tapbuf_size16_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_19_sram_inv[0:4]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size16 mux_right_track_248 (
		.in({chany_top_in[40], chany_top_in[123], chany_top_in[136], chany_top_in[232], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[52], chany_bottom_in[148], chany_bottom_in[159], chany_bottom_in[244]}),
		.sram(mux_tree_tapbuf_size16_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_20_sram_inv[0:4]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size16 mux_right_track_256 (
		.in({chany_top_in[41], chany_top_in[127], chany_top_in[137], chany_top_in[233], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[50], chany_bottom_in[146], chany_bottom_in[155], chany_bottom_in[242]}),
		.sram(mux_tree_tapbuf_size16_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_21_sram_inv[0:4]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size16 mux_right_track_264 (
		.in({chany_top_in[42], chany_top_in[131], chany_top_in[138], chany_top_in[234], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[49], chany_bottom_in[145], chany_bottom_in[151], chany_bottom_in[241]}),
		.sram(mux_tree_tapbuf_size16_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_22_sram_inv[0:4]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size16 mux_right_track_272 (
		.in({chany_top_in[44], chany_top_in[135], chany_top_in[140], chany_top_in[236], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[48], chany_bottom_in[144], chany_bottom_in[147], chany_bottom_in[240]}),
		.sram(mux_tree_tapbuf_size16_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_23_sram_inv[0:4]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size16 mux_right_track_280 (
		.in({chany_top_in[45], chany_top_in[139], chany_top_in[141], chany_top_in[237], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[46], chany_bottom_in[142:143], chany_bottom_in[238]}),
		.sram(mux_tree_tapbuf_size16_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_24_sram_inv[0:4]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size16 mux_right_track_312 (
		.in({chany_top_in[50], chany_top_in[146], chany_top_in[155], chany_top_in[242], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[41], chany_bottom_in[127], chany_bottom_in[137], chany_bottom_in[233]}),
		.sram(mux_tree_tapbuf_size16_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_25_sram_inv[0:4]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size16 mux_right_track_320 (
		.in({chany_top_in[52], chany_top_in[148], chany_top_in[159], chany_top_in[244], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[40], chany_bottom_in[123], chany_bottom_in[136], chany_bottom_in[232]}),
		.sram(mux_tree_tapbuf_size16_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_26_sram_inv[0:4]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size16 mux_right_track_328 (
		.in({chany_top_in[53], chany_top_in[149], chany_top_in[163], chany_top_in[245], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[38], chany_bottom_in[119], chany_bottom_in[134], chany_bottom_in[230]}),
		.sram(mux_tree_tapbuf_size16_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_27_sram_inv[0:4]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size16 mux_right_track_336 (
		.in({chany_top_in[54], chany_top_in[150], chany_top_in[167], chany_top_in[246], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[37], chany_bottom_in[115], chany_bottom_in[133], chany_bottom_in[229]}),
		.sram(mux_tree_tapbuf_size16_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_28_sram_inv[0:4]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size16 mux_right_track_344 (
		.in({chany_top_in[56], chany_top_in[152], chany_top_in[171], chany_top_in[248], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[36], chany_bottom_in[111], chany_bottom_in[132], chany_bottom_in[228]}),
		.sram(mux_tree_tapbuf_size16_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_29_sram_inv[0:4]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size16 mux_right_track_352 (
		.in({chany_top_in[57], chany_top_in[153], chany_top_in[175], chany_top_in[249], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[34], chany_bottom_in[107], chany_bottom_in[130], chany_bottom_in[226]}),
		.sram(mux_tree_tapbuf_size16_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_30_sram_inv[0:4]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size16 mux_right_track_384 (
		.in({chany_top_in[62], chany_top_in[158], chany_top_in[191], chany_top_in[254], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[125], chany_bottom_in[221]}),
		.sram(mux_tree_tapbuf_size16_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_31_sram_inv[0:4]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size16 mux_right_track_392 (
		.in({chany_top_in[64], chany_top_in[160], chany_top_in[195], chany_top_in[256], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[124], chany_bottom_in[220]}),
		.sram(mux_tree_tapbuf_size16_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_32_sram_inv[0:4]),
		.out(chanx_right_out[196]));

	mux_tree_tapbuf_size16 mux_right_track_400 (
		.in({chany_top_in[65], chany_top_in[161], chany_top_in[199], chany_top_in[257], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[122], chany_bottom_in[218]}),
		.sram(mux_tree_tapbuf_size16_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_33_sram_inv[0:4]),
		.out(chanx_right_out[200]));

	mux_tree_tapbuf_size16 mux_right_track_408 (
		.in({chany_top_in[66], chany_top_in[162], chany_top_in[203], chany_top_in[258], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[121], chany_bottom_in[217]}),
		.sram(mux_tree_tapbuf_size16_34_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_34_sram_inv[0:4]),
		.out(chanx_right_out[204]));

	mux_tree_tapbuf_size16 mux_right_track_416 (
		.in({chany_top_in[68], chany_top_in[164], chany_top_in[207], chany_top_in[260], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[120], chany_bottom_in[216]}),
		.sram(mux_tree_tapbuf_size16_35_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_35_sram_inv[0:4]),
		.out(chanx_right_out[208]));

	mux_tree_tapbuf_size16 mux_right_track_424 (
		.in({chany_top_in[69], chany_top_in[165], chany_top_in[211], chany_top_in[261], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[118], chany_bottom_in[214]}),
		.sram(mux_tree_tapbuf_size16_36_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_36_sram_inv[0:4]),
		.out(chanx_right_out[212]));

	mux_tree_tapbuf_size16 mux_right_track_456 (
		.in({chany_top_in[74], chany_top_in[170], chany_top_in[227], chany_top_in[266], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[113], chany_bottom_in[209]}),
		.sram(mux_tree_tapbuf_size16_37_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_37_sram_inv[0:4]),
		.out(chanx_right_out[228]));

	mux_tree_tapbuf_size16 mux_right_track_464 (
		.in({chany_top_in[76], chany_top_in[172], chany_top_in[231], chany_top_in[268], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[112], chany_bottom_in[208]}),
		.sram(mux_tree_tapbuf_size16_38_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_38_sram_inv[0:4]),
		.out(chanx_right_out[232]));

	mux_tree_tapbuf_size16 mux_right_track_472 (
		.in({chany_top_in[77], chany_top_in[173], chany_top_in[235], chany_top_in[269], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[110], chany_bottom_in[206]}),
		.sram(mux_tree_tapbuf_size16_39_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_39_sram_inv[0:4]),
		.out(chanx_right_out[236]));

	mux_tree_tapbuf_size16 mux_right_track_480 (
		.in({chany_top_in[78], chany_top_in[174], chany_top_in[239], chany_top_in[270], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[109], chany_bottom_in[205]}),
		.sram(mux_tree_tapbuf_size16_40_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_40_sram_inv[0:4]),
		.out(chanx_right_out[240]));

	mux_tree_tapbuf_size16 mux_right_track_488 (
		.in({chany_top_in[80], chany_top_in[176], chany_top_in[243], chany_top_in[272], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_42_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_51_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_69_, chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[108], chany_bottom_in[204]}),
		.sram(mux_tree_tapbuf_size16_41_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_41_sram_inv[0:4]),
		.out(chanx_right_out[244]));

	mux_tree_tapbuf_size16 mux_right_track_496 (
		.in({chany_top_in[81], chany_top_in[177], chany_top_in[247], chany_top_in[273], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[106], chany_bottom_in[202]}),
		.sram(mux_tree_tapbuf_size16_42_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_42_sram_inv[0:4]),
		.out(chanx_right_out[248]));

	mux_tree_tapbuf_size16 mux_right_track_528 (
		.in({chany_top_in[86], chany_top_in[182], chany_top_in[263], chany_top_in[278], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_38_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_47_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_65_, chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[101], chany_bottom_in[197]}),
		.sram(mux_tree_tapbuf_size16_43_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_43_sram_inv[0:4]),
		.out(chanx_right_out[264]));

	mux_tree_tapbuf_size16 mux_right_track_536 (
		.in({chany_top_in[88], chany_top_in[184], chany_top_in[267], chany_top_in[280], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_39_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_57_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_66_, chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[100], chany_bottom_in[196]}),
		.sram(mux_tree_tapbuf_size16_44_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_44_sram_inv[0:4]),
		.out(chanx_right_out[268]));

	mux_tree_tapbuf_size16 mux_right_track_544 (
		.in({chany_top_in[89], chany_top_in[185], chany_top_in[271], chany_top_in[281], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_49_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_58_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_67_, chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[98], chany_bottom_in[194]}),
		.sram(mux_tree_tapbuf_size16_45_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_45_sram_inv[0:4]),
		.out(chanx_right_out[272]));

	mux_tree_tapbuf_size16 mux_right_track_552 (
		.in({chany_top_in[90], chany_top_in[186], chany_top_in[275], chany_top_in[282], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_41_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_50_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_59_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_68_, chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[97], chany_bottom_in[193]}),
		.sram(mux_tree_tapbuf_size16_46_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_46_sram_inv[0:4]),
		.out(chanx_right_out[276]));

	mux_tree_tapbuf_size16_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_0_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_1_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_2_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_3_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_4_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_5_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_6_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_7_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_8_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_9_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_10_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_11_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_12_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_13_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_14_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_15_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_16_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_17_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_18_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_19_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_20_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_21_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_22_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_23_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_24_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_25_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_26_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_27_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_28_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_29_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_30_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_31_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_32_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_33_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_34_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_34_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_35_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_35_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_36_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_36_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_37_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_37_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_38_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_38_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_39_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_39_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_40_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_40_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_41_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_41_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_42_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_42_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_43_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_43_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_44_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_44_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_45_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_45_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_right_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_46_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_46_sram_inv[0:4]));

	mux_tree_tapbuf_size17 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[97], chany_top_in[193], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[90], chany_bottom_in[186], chany_bottom_in[275], chany_bottom_in[282]}),
		.sram(mux_tree_tapbuf_size17_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_0_sram_inv[0:4]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size17 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[106], chany_top_in[202], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[81], chany_bottom_in[177], chany_bottom_in[247], chany_bottom_in[273]}),
		.sram(mux_tree_tapbuf_size17_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_1_sram_inv[0:4]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size17 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[108], chany_top_in[204], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[80], chany_bottom_in[176], chany_bottom_in[243], chany_bottom_in[272]}),
		.sram(mux_tree_tapbuf_size17_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_2_sram_inv[0:4]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size17 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[109], chany_top_in[205], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[78], chany_bottom_in[174], chany_bottom_in[239], chany_bottom_in[270]}),
		.sram(mux_tree_tapbuf_size17_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_3_sram_inv[0:4]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size17 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[118], chany_top_in[214], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[69], chany_bottom_in[165], chany_bottom_in[211], chany_bottom_in[261]}),
		.sram(mux_tree_tapbuf_size17_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_4_sram_inv[0:4]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size17 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[120], chany_top_in[216], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[68], chany_bottom_in[164], chany_bottom_in[207], chany_bottom_in[260]}),
		.sram(mux_tree_tapbuf_size17_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_5_sram_inv[0:4]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size17 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[121], chany_top_in[217], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[66], chany_bottom_in[162], chany_bottom_in[203], chany_bottom_in[258]}),
		.sram(mux_tree_tapbuf_size17_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_6_sram_inv[0:4]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size17 mux_right_track_216 (
		.in({chany_top_in[34], chany_top_in[107], chany_top_in[130], chany_top_in[226], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[57], chany_bottom_in[153], chany_bottom_in[175], chany_bottom_in[249]}),
		.sram(mux_tree_tapbuf_size17_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_7_sram_inv[0:4]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size17 mux_right_track_224 (
		.in({chany_top_in[36], chany_top_in[111], chany_top_in[132], chany_top_in[228], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[56], chany_bottom_in[152], chany_bottom_in[171], chany_bottom_in[248]}),
		.sram(mux_tree_tapbuf_size17_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_8_sram_inv[0:4]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size17 mux_right_track_232 (
		.in({chany_top_in[37], chany_top_in[115], chany_top_in[133], chany_top_in[229], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[54], chany_bottom_in[150], chany_bottom_in[167], chany_bottom_in[246]}),
		.sram(mux_tree_tapbuf_size17_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_9_sram_inv[0:4]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size17 mux_right_track_288 (
		.in({chany_top_in[46], chany_top_in[142:143], chany_top_in[238], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[45], chany_bottom_in[139], chany_bottom_in[141], chany_bottom_in[237]}),
		.sram(mux_tree_tapbuf_size17_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_10_sram_inv[0:4]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size17 mux_right_track_296 (
		.in({chany_top_in[48], chany_top_in[144], chany_top_in[147], chany_top_in[240], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[44], chany_bottom_in[135], chany_bottom_in[140], chany_bottom_in[236]}),
		.sram(mux_tree_tapbuf_size17_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_11_sram_inv[0:4]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size17 mux_right_track_304 (
		.in({chany_top_in[49], chany_top_in[145], chany_top_in[151], chany_top_in[241], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[42], chany_bottom_in[131], chany_bottom_in[138], chany_bottom_in[234]}),
		.sram(mux_tree_tapbuf_size17_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_12_sram_inv[0:4]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size17 mux_right_track_360 (
		.in({chany_top_in[58], chany_top_in[154], chany_top_in[179], chany_top_in[250], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[33], chany_bottom_in[103], chany_bottom_in[129], chany_bottom_in[225]}),
		.sram(mux_tree_tapbuf_size17_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_13_sram_inv[0:4]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size17 mux_right_track_368 (
		.in({chany_top_in[60], chany_top_in[156], chany_top_in[183], chany_top_in[252], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[32], chany_bottom_in[99], chany_bottom_in[128], chany_bottom_in[224]}),
		.sram(mux_tree_tapbuf_size17_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_14_sram_inv[0:4]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size17 mux_right_track_376 (
		.in({chany_top_in[61], chany_top_in[157], chany_top_in[187], chany_top_in[253], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[30], chany_bottom_in[95], chany_bottom_in[126], chany_bottom_in[222]}),
		.sram(mux_tree_tapbuf_size17_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_15_sram_inv[0:4]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size17 mux_right_track_432 (
		.in({chany_top_in[70], chany_top_in[166], chany_top_in[215], chany_top_in[262], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[117], chany_bottom_in[213]}),
		.sram(mux_tree_tapbuf_size17_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_16_sram_inv[0:4]),
		.out(chanx_right_out[216]));

	mux_tree_tapbuf_size17 mux_right_track_440 (
		.in({chany_top_in[72], chany_top_in[168], chany_top_in[219], chany_top_in[264], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[116], chany_bottom_in[212]}),
		.sram(mux_tree_tapbuf_size17_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_17_sram_inv[0:4]),
		.out(chanx_right_out[220]));

	mux_tree_tapbuf_size17 mux_right_track_448 (
		.in({chany_top_in[73], chany_top_in[169], chany_top_in[223], chany_top_in[265], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[114], chany_bottom_in[210]}),
		.sram(mux_tree_tapbuf_size17_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_18_sram_inv[0:4]),
		.out(chanx_right_out[224]));

	mux_tree_tapbuf_size17 mux_right_track_504 (
		.in({chany_top_in[82], chany_top_in[178], chany_top_in[251], chany_top_in[274], right_top_grid_bottom_width_0_height_0_subtile_0__pin_error_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_35_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_53_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_62_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_1_, chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[105], chany_bottom_in[201]}),
		.sram(mux_tree_tapbuf_size17_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_19_sram_inv[0:4]),
		.out(chanx_right_out[252]));

	mux_tree_tapbuf_size17 mux_right_track_512 (
		.in({chany_top_in[84], chany_top_in[180], chany_top_in[255], chany_top_in[276], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_45_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_54_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_63_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_2_, chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[104], chany_bottom_in[200]}),
		.sram(mux_tree_tapbuf_size17_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_20_sram_inv[0:4]),
		.out(chanx_right_out[256]));

	mux_tree_tapbuf_size17 mux_right_track_520 (
		.in({chany_top_in[85], chany_top_in[181], chany_top_in[259], chany_top_in[277], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_37_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_46_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_55_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_64_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[102], chany_bottom_in[198]}),
		.sram(mux_tree_tapbuf_size17_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_21_sram_inv[0:4]),
		.out(chanx_right_out[260]));

	mux_tree_tapbuf_size17_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_0_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_1_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_2_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_3_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_4_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_5_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_6_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_7_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_8_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_9_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_10_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_11_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_12_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_13_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_14_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_15_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_16_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_17_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_18_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_19_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_20_sram_inv[0:4]));

	mux_tree_tapbuf_size17_mem mem_right_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_21_sram_inv[0:4]));

	mux_tree_tapbuf_size14 mux_right_track_568 (
		.in({chany_top_in[93], chany_top_in[189], chany_top_in[283], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_43_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_2_61_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_0_, chany_bottom_in[94], chany_bottom_in[190], chany_bottom_in[284]}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chanx_right_out[284]));

	mux_tree_tapbuf_size14_mem mem_right_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size8 mux_bottom_track_1 (
		.in({chanx_right_in[93], chanx_right_in[189], chanx_right_in[283], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[1], chanx_left_in[7], chanx_left_in[97], chanx_left_in[193]}),
		.sram(mux_tree_tapbuf_size8_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_0_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size8 mux_bottom_track_9 (
		.in({chanx_right_in[92], chanx_right_in[188], chanx_right_in[279], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[2], chanx_left_in[11], chanx_left_in[98], chanx_left_in[194]}),
		.sram(mux_tree_tapbuf_size8_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_1_sram_inv[0:3]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size8 mux_bottom_track_17 (
		.in({chanx_right_in[90], chanx_right_in[186], chanx_right_in[275], chanx_right_in[282], chanx_left_in[4], chanx_left_in[15], chanx_left_in[100], chanx_left_in[196]}),
		.sram(mux_tree_tapbuf_size8_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_2_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size8 mux_bottom_track_25 (
		.in({chanx_right_in[89], chanx_right_in[185], chanx_right_in[271], chanx_right_in[281], chanx_left_in[5], chanx_left_in[19], chanx_left_in[101], chanx_left_in[197]}),
		.sram(mux_tree_tapbuf_size8_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_3_sram_inv[0:3]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size8 mux_bottom_track_33 (
		.in({chanx_right_in[88], chanx_right_in[184], chanx_right_in[267], chanx_right_in[280], chanx_left_in[6], chanx_left_in[23], chanx_left_in[102], chanx_left_in[198]}),
		.sram(mux_tree_tapbuf_size8_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_4_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size8 mux_bottom_track_41 (
		.in({chanx_right_in[86], chanx_right_in[182], chanx_right_in[263], chanx_right_in[278], chanx_left_in[8], chanx_left_in[27], chanx_left_in[104], chanx_left_in[200]}),
		.sram(mux_tree_tapbuf_size8_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_5_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size8 mux_bottom_track_49 (
		.in({chanx_right_in[85], chanx_right_in[181], chanx_right_in[259], chanx_right_in[277], chanx_left_in[9], chanx_left_in[31], chanx_left_in[105], chanx_left_in[201]}),
		.sram(mux_tree_tapbuf_size8_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_6_sram_inv[0:3]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size8 mux_bottom_track_57 (
		.in({chanx_right_in[84], chanx_right_in[180], chanx_right_in[255], chanx_right_in[276], chanx_left_in[10], chanx_left_in[35], chanx_left_in[106], chanx_left_in[202]}),
		.sram(mux_tree_tapbuf_size8_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_7_sram_inv[0:3]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size8 mux_bottom_track_65 (
		.in({chanx_right_in[82], chanx_right_in[178], chanx_right_in[251], chanx_right_in[274], chanx_left_in[12], chanx_left_in[39], chanx_left_in[108], chanx_left_in[204]}),
		.sram(mux_tree_tapbuf_size8_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_8_sram_inv[0:3]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size8 mux_bottom_track_89 (
		.in({chanx_right_in[78], chanx_right_in[174], chanx_right_in[239], chanx_right_in[270], chanx_left_in[16], chanx_left_in[51], chanx_left_in[112], chanx_left_in[208]}),
		.sram(mux_tree_tapbuf_size8_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_9_sram_inv[0:3]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size8 mux_bottom_track_97 (
		.in({chanx_right_in[77], chanx_right_in[173], chanx_right_in[235], chanx_right_in[269], chanx_left_in[17], chanx_left_in[55], chanx_left_in[113], chanx_left_in[209]}),
		.sram(mux_tree_tapbuf_size8_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_10_sram_inv[0:3]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size8 mux_bottom_track_105 (
		.in({chanx_right_in[76], chanx_right_in[172], chanx_right_in[231], chanx_right_in[268], chanx_left_in[18], chanx_left_in[59], chanx_left_in[114], chanx_left_in[210]}),
		.sram(mux_tree_tapbuf_size8_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_11_sram_inv[0:3]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size8 mux_bottom_track_113 (
		.in({chanx_right_in[74], chanx_right_in[170], chanx_right_in[227], chanx_right_in[266], chanx_left_in[20], chanx_left_in[63], chanx_left_in[116], chanx_left_in[212]}),
		.sram(mux_tree_tapbuf_size8_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_12_sram_inv[0:3]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size8 mux_bottom_track_121 (
		.in({chanx_right_in[73], chanx_right_in[169], chanx_right_in[223], chanx_right_in[265], chanx_left_in[21], chanx_left_in[67], chanx_left_in[117], chanx_left_in[213]}),
		.sram(mux_tree_tapbuf_size8_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_13_sram_inv[0:3]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size8 mux_bottom_track_129 (
		.in({chanx_right_in[72], chanx_right_in[168], chanx_right_in[219], chanx_right_in[264], chanx_left_in[22], chanx_left_in[71], chanx_left_in[118], chanx_left_in[214]}),
		.sram(mux_tree_tapbuf_size8_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_14_sram_inv[0:3]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size8 mux_bottom_track_137 (
		.in({chanx_right_in[70], chanx_right_in[166], chanx_right_in[215], chanx_right_in[262], chanx_left_in[24], chanx_left_in[75], chanx_left_in[120], chanx_left_in[216]}),
		.sram(mux_tree_tapbuf_size8_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_15_sram_inv[0:3]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size8 mux_bottom_track_161 (
		.in({chanx_right_in[66], chanx_right_in[162], chanx_right_in[203], chanx_right_in[258], chanx_left_in[28], chanx_left_in[87], chanx_left_in[124], chanx_left_in[220]}),
		.sram(mux_tree_tapbuf_size8_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_16_sram_inv[0:3]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size8 mux_bottom_track_169 (
		.in({chanx_right_in[65], chanx_right_in[161], chanx_right_in[199], chanx_right_in[257], chanx_left_in[29], chanx_left_in[91], chanx_left_in[125], chanx_left_in[221]}),
		.sram(mux_tree_tapbuf_size8_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_17_sram_inv[0:3]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size8 mux_bottom_track_177 (
		.in({chanx_right_in[64], chanx_right_in[160], chanx_right_in[195], chanx_right_in[256], chanx_left_in[30], chanx_left_in[95], chanx_left_in[126], chanx_left_in[222]}),
		.sram(mux_tree_tapbuf_size8_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_18_sram_inv[0:3]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size8 mux_bottom_track_185 (
		.in({chanx_right_in[62], chanx_right_in[158], chanx_right_in[191], chanx_right_in[254], chanx_left_in[32], chanx_left_in[99], chanx_left_in[128], chanx_left_in[224]}),
		.sram(mux_tree_tapbuf_size8_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_19_sram_inv[0:3]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size8 mux_bottom_track_193 (
		.in({chanx_right_in[61], chanx_right_in[157], chanx_right_in[187], chanx_right_in[253], chanx_left_in[33], chanx_left_in[103], chanx_left_in[129], chanx_left_in[225]}),
		.sram(mux_tree_tapbuf_size8_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_20_sram_inv[0:3]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size8 mux_bottom_track_201 (
		.in({chanx_right_in[60], chanx_right_in[156], chanx_right_in[183], chanx_right_in[252], chanx_left_in[34], chanx_left_in[107], chanx_left_in[130], chanx_left_in[226]}),
		.sram(mux_tree_tapbuf_size8_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_21_sram_inv[0:3]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size8 mux_bottom_track_209 (
		.in({chanx_right_in[58], chanx_right_in[154], chanx_right_in[179], chanx_right_in[250], chanx_left_in[36], chanx_left_in[111], chanx_left_in[132], chanx_left_in[228]}),
		.sram(mux_tree_tapbuf_size8_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_22_sram_inv[0:3]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size8 mux_bottom_track_233 (
		.in({chanx_right_in[54], chanx_right_in[150], chanx_right_in[167], chanx_right_in[246], chanx_left_in[40], chanx_left_in[123], chanx_left_in[136], chanx_left_in[232]}),
		.sram(mux_tree_tapbuf_size8_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_23_sram_inv[0:3]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size8 mux_bottom_track_241 (
		.in({chanx_right_in[53], chanx_right_in[149], chanx_right_in[163], chanx_right_in[245], chanx_left_in[41], chanx_left_in[127], chanx_left_in[137], chanx_left_in[233]}),
		.sram(mux_tree_tapbuf_size8_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_24_sram_inv[0:3]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size8 mux_bottom_track_249 (
		.in({chanx_right_in[52], chanx_right_in[148], chanx_right_in[159], chanx_right_in[244], chanx_left_in[42], chanx_left_in[131], chanx_left_in[138], chanx_left_in[234]}),
		.sram(mux_tree_tapbuf_size8_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_25_sram_inv[0:3]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size8 mux_bottom_track_257 (
		.in({chanx_right_in[50], chanx_right_in[146], chanx_right_in[155], chanx_right_in[242], chanx_left_in[44], chanx_left_in[135], chanx_left_in[140], chanx_left_in[236]}),
		.sram(mux_tree_tapbuf_size8_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_26_sram_inv[0:3]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size8 mux_bottom_track_265 (
		.in({chanx_right_in[49], chanx_right_in[145], chanx_right_in[151], chanx_right_in[241], chanx_left_in[45], chanx_left_in[139], chanx_left_in[141], chanx_left_in[237]}),
		.sram(mux_tree_tapbuf_size8_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_27_sram_inv[0:3]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size8 mux_bottom_track_273 (
		.in({chanx_right_in[48], chanx_right_in[144], chanx_right_in[147], chanx_right_in[240], chanx_left_in[46], chanx_left_in[142:143], chanx_left_in[238]}),
		.sram(mux_tree_tapbuf_size8_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_28_sram_inv[0:3]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size8 mux_bottom_track_281 (
		.in({chanx_right_in[46], chanx_right_in[142:143], chanx_right_in[238], chanx_left_in[48], chanx_left_in[144], chanx_left_in[147], chanx_left_in[240]}),
		.sram(mux_tree_tapbuf_size8_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_29_sram_inv[0:3]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size8 mux_bottom_track_305 (
		.in({chanx_right_in[42], chanx_right_in[131], chanx_right_in[138], chanx_right_in[234], chanx_left_in[52], chanx_left_in[148], chanx_left_in[159], chanx_left_in[244]}),
		.sram(mux_tree_tapbuf_size8_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_30_sram_inv[0:3]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size8 mux_bottom_track_313 (
		.in({chanx_right_in[41], chanx_right_in[127], chanx_right_in[137], chanx_right_in[233], chanx_left_in[53], chanx_left_in[149], chanx_left_in[163], chanx_left_in[245]}),
		.sram(mux_tree_tapbuf_size8_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_31_sram_inv[0:3]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size8 mux_bottom_track_321 (
		.in({chanx_right_in[40], chanx_right_in[123], chanx_right_in[136], chanx_right_in[232], chanx_left_in[54], chanx_left_in[150], chanx_left_in[167], chanx_left_in[246]}),
		.sram(mux_tree_tapbuf_size8_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_32_sram_inv[0:3]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size8 mux_bottom_track_329 (
		.in({chanx_right_in[38], chanx_right_in[119], chanx_right_in[134], chanx_right_in[230], chanx_left_in[56], chanx_left_in[152], chanx_left_in[171], chanx_left_in[248]}),
		.sram(mux_tree_tapbuf_size8_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_33_sram_inv[0:3]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size8 mux_bottom_track_337 (
		.in({chanx_right_in[37], chanx_right_in[115], chanx_right_in[133], chanx_right_in[229], chanx_left_in[57], chanx_left_in[153], chanx_left_in[175], chanx_left_in[249]}),
		.sram(mux_tree_tapbuf_size8_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_34_sram_inv[0:3]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size8 mux_bottom_track_345 (
		.in({chanx_right_in[36], chanx_right_in[111], chanx_right_in[132], chanx_right_in[228], chanx_left_in[58], chanx_left_in[154], chanx_left_in[179], chanx_left_in[250]}),
		.sram(mux_tree_tapbuf_size8_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_35_sram_inv[0:3]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size8 mux_bottom_track_353 (
		.in({chanx_right_in[34], chanx_right_in[107], chanx_right_in[130], chanx_right_in[226], chanx_left_in[60], chanx_left_in[156], chanx_left_in[183], chanx_left_in[252]}),
		.sram(mux_tree_tapbuf_size8_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_36_sram_inv[0:3]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size8 mux_bottom_track_377 (
		.in({chanx_right_in[30], chanx_right_in[95], chanx_right_in[126], chanx_right_in[222], chanx_left_in[64], chanx_left_in[160], chanx_left_in[195], chanx_left_in[256]}),
		.sram(mux_tree_tapbuf_size8_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_37_sram_inv[0:3]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size8 mux_bottom_track_385 (
		.in({chanx_right_in[29], chanx_right_in[91], chanx_right_in[125], chanx_right_in[221], chanx_left_in[65], chanx_left_in[161], chanx_left_in[199], chanx_left_in[257]}),
		.sram(mux_tree_tapbuf_size8_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_38_sram_inv[0:3]),
		.out(chany_bottom_out[192]));

	mux_tree_tapbuf_size8 mux_bottom_track_393 (
		.in({chanx_right_in[28], chanx_right_in[87], chanx_right_in[124], chanx_right_in[220], chanx_left_in[66], chanx_left_in[162], chanx_left_in[203], chanx_left_in[258]}),
		.sram(mux_tree_tapbuf_size8_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_39_sram_inv[0:3]),
		.out(chany_bottom_out[196]));

	mux_tree_tapbuf_size8 mux_bottom_track_401 (
		.in({chanx_right_in[26], chanx_right_in[83], chanx_right_in[122], chanx_right_in[218], chanx_left_in[68], chanx_left_in[164], chanx_left_in[207], chanx_left_in[260]}),
		.sram(mux_tree_tapbuf_size8_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_40_sram_inv[0:3]),
		.out(chany_bottom_out[200]));

	mux_tree_tapbuf_size8 mux_bottom_track_409 (
		.in({chanx_right_in[25], chanx_right_in[79], chanx_right_in[121], chanx_right_in[217], chanx_left_in[69], chanx_left_in[165], chanx_left_in[211], chanx_left_in[261]}),
		.sram(mux_tree_tapbuf_size8_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_41_sram_inv[0:3]),
		.out(chany_bottom_out[204]));

	mux_tree_tapbuf_size8 mux_bottom_track_417 (
		.in({chanx_right_in[24], chanx_right_in[75], chanx_right_in[120], chanx_right_in[216], chanx_left_in[70], chanx_left_in[166], chanx_left_in[215], chanx_left_in[262]}),
		.sram(mux_tree_tapbuf_size8_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_42_sram_inv[0:3]),
		.out(chany_bottom_out[208]));

	mux_tree_tapbuf_size8 mux_bottom_track_425 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[118], chanx_right_in[214], chanx_left_in[72], chanx_left_in[168], chanx_left_in[219], chanx_left_in[264]}),
		.sram(mux_tree_tapbuf_size8_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_43_sram_inv[0:3]),
		.out(chany_bottom_out[212]));

	mux_tree_tapbuf_size8 mux_bottom_track_449 (
		.in({chanx_right_in[18], chanx_right_in[59], chanx_right_in[114], chanx_right_in[210], chanx_left_in[76], chanx_left_in[172], chanx_left_in[231], chanx_left_in[268]}),
		.sram(mux_tree_tapbuf_size8_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_44_sram_inv[0:3]),
		.out(chany_bottom_out[224]));

	mux_tree_tapbuf_size8 mux_bottom_track_457 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[113], chanx_right_in[209], chanx_left_in[77], chanx_left_in[173], chanx_left_in[235], chanx_left_in[269]}),
		.sram(mux_tree_tapbuf_size8_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_45_sram_inv[0:3]),
		.out(chany_bottom_out[228]));

	mux_tree_tapbuf_size8 mux_bottom_track_465 (
		.in({chanx_right_in[16], chanx_right_in[51], chanx_right_in[112], chanx_right_in[208], chanx_left_in[78], chanx_left_in[174], chanx_left_in[239], chanx_left_in[270]}),
		.sram(mux_tree_tapbuf_size8_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_46_sram_inv[0:3]),
		.out(chany_bottom_out[232]));

	mux_tree_tapbuf_size8 mux_bottom_track_473 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[110], chanx_right_in[206], chanx_left_in[80], chanx_left_in[176], chanx_left_in[243], chanx_left_in[272]}),
		.sram(mux_tree_tapbuf_size8_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_47_sram_inv[0:3]),
		.out(chany_bottom_out[236]));

	mux_tree_tapbuf_size8 mux_bottom_track_481 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[109], chanx_right_in[205], chanx_left_in[81], chanx_left_in[177], chanx_left_in[247], chanx_left_in[273]}),
		.sram(mux_tree_tapbuf_size8_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_48_sram_inv[0:3]),
		.out(chany_bottom_out[240]));

	mux_tree_tapbuf_size8 mux_bottom_track_489 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[108], chanx_right_in[204], chanx_left_in[82], chanx_left_in[178], chanx_left_in[251], chanx_left_in[274]}),
		.sram(mux_tree_tapbuf_size8_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_49_sram_inv[0:3]),
		.out(chany_bottom_out[244]));

	mux_tree_tapbuf_size8 mux_bottom_track_497 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[106], chanx_right_in[202], chanx_left_in[84], chanx_left_in[180], chanx_left_in[255], chanx_left_in[276]}),
		.sram(mux_tree_tapbuf_size8_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_50_sram_inv[0:3]),
		.out(chany_bottom_out[248]));

	mux_tree_tapbuf_size8 mux_bottom_track_521 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[102], chanx_right_in[198], chanx_left_in[88], chanx_left_in[184], chanx_left_in[267], chanx_left_in[280]}),
		.sram(mux_tree_tapbuf_size8_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_51_sram_inv[0:3]),
		.out(chany_bottom_out[260]));

	mux_tree_tapbuf_size8 mux_bottom_track_529 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[101], chanx_right_in[197], chanx_left_in[89], chanx_left_in[185], chanx_left_in[271], chanx_left_in[281]}),
		.sram(mux_tree_tapbuf_size8_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_52_sram_inv[0:3]),
		.out(chany_bottom_out[264]));

	mux_tree_tapbuf_size8 mux_bottom_track_537 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[100], chanx_right_in[196], chanx_left_in[90], chanx_left_in[186], chanx_left_in[275], chanx_left_in[282]}),
		.sram(mux_tree_tapbuf_size8_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_53_sram_inv[0:3]),
		.out(chany_bottom_out[268]));

	mux_tree_tapbuf_size8 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[96], chany_top_in[192], chany_bottom_in[94], chany_bottom_in[190], chany_bottom_in[284], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size8_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_54_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size8 mux_left_track_9 (
		.in({chany_top_in[94], chany_top_in[190], chany_top_in[284], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[96], chany_bottom_in[192], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size8_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_55_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size8 mux_left_track_33 (
		.in({chany_top_in[90], chany_top_in[186], chany_top_in[275], chany_top_in[282], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[100], chany_bottom_in[196]}),
		.sram(mux_tree_tapbuf_size8_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_56_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size8 mux_left_track_41 (
		.in({chany_top_in[89], chany_top_in[185], chany_top_in[271], chany_top_in[281], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[101], chany_bottom_in[197]}),
		.sram(mux_tree_tapbuf_size8_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_57_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size8 mux_left_track_49 (
		.in({chany_top_in[88], chany_top_in[184], chany_top_in[267], chany_top_in[280], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[102], chany_bottom_in[198]}),
		.sram(mux_tree_tapbuf_size8_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_58_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size8 mux_left_track_57 (
		.in({chany_top_in[86], chany_top_in[182], chany_top_in[263], chany_top_in[278], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[104], chany_bottom_in[200]}),
		.sram(mux_tree_tapbuf_size8_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_59_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size8 mux_left_track_65 (
		.in({chany_top_in[85], chany_top_in[181], chany_top_in[259], chany_top_in[277], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[105], chany_bottom_in[201]}),
		.sram(mux_tree_tapbuf_size8_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_60_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size8 mux_left_track_89 (
		.in({chany_top_in[81], chany_top_in[177], chany_top_in[247], chany_top_in[273], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[109], chany_bottom_in[205]}),
		.sram(mux_tree_tapbuf_size8_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_61_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size8 mux_left_track_97 (
		.in({chany_top_in[80], chany_top_in[176], chany_top_in[243], chany_top_in[272], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[110], chany_bottom_in[206]}),
		.sram(mux_tree_tapbuf_size8_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_62_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size8 mux_left_track_105 (
		.in({chany_top_in[78], chany_top_in[174], chany_top_in[239], chany_top_in[270], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[112], chany_bottom_in[208]}),
		.sram(mux_tree_tapbuf_size8_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_63_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size8 mux_left_track_113 (
		.in({chany_top_in[77], chany_top_in[173], chany_top_in[235], chany_top_in[269], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[113], chany_bottom_in[209]}),
		.sram(mux_tree_tapbuf_size8_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_64_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size8 mux_left_track_121 (
		.in({chany_top_in[76], chany_top_in[172], chany_top_in[231], chany_top_in[268], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[114], chany_bottom_in[210]}),
		.sram(mux_tree_tapbuf_size8_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_65_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size8 mux_left_track_129 (
		.in({chany_top_in[74], chany_top_in[170], chany_top_in[227], chany_top_in[266], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[116], chany_bottom_in[212]}),
		.sram(mux_tree_tapbuf_size8_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_66_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size8 mux_left_track_137 (
		.in({chany_top_in[73], chany_top_in[169], chany_top_in[223], chany_top_in[265], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[117], chany_bottom_in[213]}),
		.sram(mux_tree_tapbuf_size8_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_67_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size8 mux_left_track_161 (
		.in({chany_top_in[69], chany_top_in[165], chany_top_in[211], chany_top_in[261], chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[121], chany_bottom_in[217]}),
		.sram(mux_tree_tapbuf_size8_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_68_sram_inv[0:3]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size8 mux_left_track_169 (
		.in({chany_top_in[68], chany_top_in[164], chany_top_in[207], chany_top_in[260], chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[122], chany_bottom_in[218]}),
		.sram(mux_tree_tapbuf_size8_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_69_sram_inv[0:3]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size8 mux_left_track_177 (
		.in({chany_top_in[66], chany_top_in[162], chany_top_in[203], chany_top_in[258], chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[124], chany_bottom_in[220]}),
		.sram(mux_tree_tapbuf_size8_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_70_sram_inv[0:3]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size8 mux_left_track_185 (
		.in({chany_top_in[65], chany_top_in[161], chany_top_in[199], chany_top_in[257], chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[125], chany_bottom_in[221]}),
		.sram(mux_tree_tapbuf_size8_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_71_sram_inv[0:3]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size8 mux_left_track_193 (
		.in({chany_top_in[64], chany_top_in[160], chany_top_in[195], chany_top_in[256], chany_bottom_in[30], chany_bottom_in[95], chany_bottom_in[126], chany_bottom_in[222]}),
		.sram(mux_tree_tapbuf_size8_72_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_72_sram_inv[0:3]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size8 mux_left_track_201 (
		.in({chany_top_in[62], chany_top_in[158], chany_top_in[191], chany_top_in[254], chany_bottom_in[32], chany_bottom_in[99], chany_bottom_in[128], chany_bottom_in[224]}),
		.sram(mux_tree_tapbuf_size8_73_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_73_sram_inv[0:3]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size8 mux_left_track_209 (
		.in({chany_top_in[61], chany_top_in[157], chany_top_in[187], chany_top_in[253], chany_bottom_in[33], chany_bottom_in[103], chany_bottom_in[129], chany_bottom_in[225]}),
		.sram(mux_tree_tapbuf_size8_74_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_74_sram_inv[0:3]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size8 mux_left_track_233 (
		.in({chany_top_in[57], chany_top_in[153], chany_top_in[175], chany_top_in[249], chany_bottom_in[37], chany_bottom_in[115], chany_bottom_in[133], chany_bottom_in[229]}),
		.sram(mux_tree_tapbuf_size8_75_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_75_sram_inv[0:3]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size8 mux_left_track_241 (
		.in({chany_top_in[56], chany_top_in[152], chany_top_in[171], chany_top_in[248], chany_bottom_in[38], chany_bottom_in[119], chany_bottom_in[134], chany_bottom_in[230]}),
		.sram(mux_tree_tapbuf_size8_76_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_76_sram_inv[0:3]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size8 mux_left_track_249 (
		.in({chany_top_in[54], chany_top_in[150], chany_top_in[167], chany_top_in[246], chany_bottom_in[40], chany_bottom_in[123], chany_bottom_in[136], chany_bottom_in[232]}),
		.sram(mux_tree_tapbuf_size8_77_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_77_sram_inv[0:3]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size8 mux_left_track_257 (
		.in({chany_top_in[53], chany_top_in[149], chany_top_in[163], chany_top_in[245], chany_bottom_in[41], chany_bottom_in[127], chany_bottom_in[137], chany_bottom_in[233]}),
		.sram(mux_tree_tapbuf_size8_78_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_78_sram_inv[0:3]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size8 mux_left_track_265 (
		.in({chany_top_in[52], chany_top_in[148], chany_top_in[159], chany_top_in[244], chany_bottom_in[42], chany_bottom_in[131], chany_bottom_in[138], chany_bottom_in[234]}),
		.sram(mux_tree_tapbuf_size8_79_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_79_sram_inv[0:3]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size8 mux_left_track_273 (
		.in({chany_top_in[50], chany_top_in[146], chany_top_in[155], chany_top_in[242], chany_bottom_in[44], chany_bottom_in[135], chany_bottom_in[140], chany_bottom_in[236]}),
		.sram(mux_tree_tapbuf_size8_80_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_80_sram_inv[0:3]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size8 mux_left_track_281 (
		.in({chany_top_in[49], chany_top_in[145], chany_top_in[151], chany_top_in[241], chany_bottom_in[45], chany_bottom_in[139], chany_bottom_in[141], chany_bottom_in[237]}),
		.sram(mux_tree_tapbuf_size8_81_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_81_sram_inv[0:3]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size8 mux_left_track_305 (
		.in({chany_top_in[45], chany_top_in[139], chany_top_in[141], chany_top_in[237], chany_bottom_in[49], chany_bottom_in[145], chany_bottom_in[151], chany_bottom_in[241]}),
		.sram(mux_tree_tapbuf_size8_82_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_82_sram_inv[0:3]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size8 mux_left_track_313 (
		.in({chany_top_in[44], chany_top_in[135], chany_top_in[140], chany_top_in[236], chany_bottom_in[50], chany_bottom_in[146], chany_bottom_in[155], chany_bottom_in[242]}),
		.sram(mux_tree_tapbuf_size8_83_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_83_sram_inv[0:3]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size8 mux_left_track_321 (
		.in({chany_top_in[42], chany_top_in[131], chany_top_in[138], chany_top_in[234], chany_bottom_in[52], chany_bottom_in[148], chany_bottom_in[159], chany_bottom_in[244]}),
		.sram(mux_tree_tapbuf_size8_84_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_84_sram_inv[0:3]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size8 mux_left_track_329 (
		.in({chany_top_in[41], chany_top_in[127], chany_top_in[137], chany_top_in[233], chany_bottom_in[53], chany_bottom_in[149], chany_bottom_in[163], chany_bottom_in[245]}),
		.sram(mux_tree_tapbuf_size8_85_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_85_sram_inv[0:3]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size8 mux_left_track_337 (
		.in({chany_top_in[40], chany_top_in[123], chany_top_in[136], chany_top_in[232], chany_bottom_in[54], chany_bottom_in[150], chany_bottom_in[167], chany_bottom_in[246]}),
		.sram(mux_tree_tapbuf_size8_86_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_86_sram_inv[0:3]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size8 mux_left_track_345 (
		.in({chany_top_in[38], chany_top_in[119], chany_top_in[134], chany_top_in[230], chany_bottom_in[56], chany_bottom_in[152], chany_bottom_in[171], chany_bottom_in[248]}),
		.sram(mux_tree_tapbuf_size8_87_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_87_sram_inv[0:3]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size8 mux_left_track_353 (
		.in({chany_top_in[37], chany_top_in[115], chany_top_in[133], chany_top_in[229], chany_bottom_in[57], chany_bottom_in[153], chany_bottom_in[175], chany_bottom_in[249]}),
		.sram(mux_tree_tapbuf_size8_88_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_88_sram_inv[0:3]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size8 mux_left_track_377 (
		.in({chany_top_in[33], chany_top_in[103], chany_top_in[129], chany_top_in[225], chany_bottom_in[61], chany_bottom_in[157], chany_bottom_in[187], chany_bottom_in[253]}),
		.sram(mux_tree_tapbuf_size8_89_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_89_sram_inv[0:3]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size8 mux_left_track_385 (
		.in({chany_top_in[32], chany_top_in[99], chany_top_in[128], chany_top_in[224], chany_bottom_in[62], chany_bottom_in[158], chany_bottom_in[191], chany_bottom_in[254]}),
		.sram(mux_tree_tapbuf_size8_90_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_90_sram_inv[0:3]),
		.out(chanx_left_out[192]));

	mux_tree_tapbuf_size8 mux_left_track_393 (
		.in({chany_top_in[30], chany_top_in[95], chany_top_in[126], chany_top_in[222], chany_bottom_in[64], chany_bottom_in[160], chany_bottom_in[195], chany_bottom_in[256]}),
		.sram(mux_tree_tapbuf_size8_91_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_91_sram_inv[0:3]),
		.out(chanx_left_out[196]));

	mux_tree_tapbuf_size8 mux_left_track_401 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[125], chany_top_in[221], chany_bottom_in[65], chany_bottom_in[161], chany_bottom_in[199], chany_bottom_in[257]}),
		.sram(mux_tree_tapbuf_size8_92_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_92_sram_inv[0:3]),
		.out(chanx_left_out[200]));

	mux_tree_tapbuf_size8 mux_left_track_409 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[124], chany_top_in[220], chany_bottom_in[66], chany_bottom_in[162], chany_bottom_in[203], chany_bottom_in[258]}),
		.sram(mux_tree_tapbuf_size8_93_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_93_sram_inv[0:3]),
		.out(chanx_left_out[204]));

	mux_tree_tapbuf_size8 mux_left_track_417 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[122], chany_top_in[218], chany_bottom_in[68], chany_bottom_in[164], chany_bottom_in[207], chany_bottom_in[260]}),
		.sram(mux_tree_tapbuf_size8_94_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_94_sram_inv[0:3]),
		.out(chanx_left_out[208]));

	mux_tree_tapbuf_size8 mux_left_track_425 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[121], chany_top_in[217], chany_bottom_in[69], chany_bottom_in[165], chany_bottom_in[211], chany_bottom_in[261]}),
		.sram(mux_tree_tapbuf_size8_95_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_95_sram_inv[0:3]),
		.out(chanx_left_out[212]));

	mux_tree_tapbuf_size8 mux_left_track_449 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[117], chany_top_in[213], chany_bottom_in[73], chany_bottom_in[169], chany_bottom_in[223], chany_bottom_in[265]}),
		.sram(mux_tree_tapbuf_size8_96_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_96_sram_inv[0:3]),
		.out(chanx_left_out[224]));

	mux_tree_tapbuf_size8 mux_left_track_457 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[116], chany_top_in[212], chany_bottom_in[74], chany_bottom_in[170], chany_bottom_in[227], chany_bottom_in[266]}),
		.sram(mux_tree_tapbuf_size8_97_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_97_sram_inv[0:3]),
		.out(chanx_left_out[228]));

	mux_tree_tapbuf_size8 mux_left_track_465 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[114], chany_top_in[210], chany_bottom_in[76], chany_bottom_in[172], chany_bottom_in[231], chany_bottom_in[268]}),
		.sram(mux_tree_tapbuf_size8_98_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_98_sram_inv[0:3]),
		.out(chanx_left_out[232]));

	mux_tree_tapbuf_size8 mux_left_track_473 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[113], chany_top_in[209], chany_bottom_in[77], chany_bottom_in[173], chany_bottom_in[235], chany_bottom_in[269]}),
		.sram(mux_tree_tapbuf_size8_99_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_99_sram_inv[0:3]),
		.out(chanx_left_out[236]));

	mux_tree_tapbuf_size8 mux_left_track_481 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[112], chany_top_in[208], chany_bottom_in[78], chany_bottom_in[174], chany_bottom_in[239], chany_bottom_in[270]}),
		.sram(mux_tree_tapbuf_size8_100_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_100_sram_inv[0:3]),
		.out(chanx_left_out[240]));

	mux_tree_tapbuf_size8 mux_left_track_489 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[110], chany_top_in[206], chany_bottom_in[80], chany_bottom_in[176], chany_bottom_in[243], chany_bottom_in[272]}),
		.sram(mux_tree_tapbuf_size8_101_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_101_sram_inv[0:3]),
		.out(chanx_left_out[244]));

	mux_tree_tapbuf_size8 mux_left_track_497 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[109], chany_top_in[205], chany_bottom_in[81], chany_bottom_in[177], chany_bottom_in[247], chany_bottom_in[273]}),
		.sram(mux_tree_tapbuf_size8_102_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_102_sram_inv[0:3]),
		.out(chanx_left_out[248]));

	mux_tree_tapbuf_size8 mux_left_track_521 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[105], chany_top_in[201], chany_bottom_in[85], chany_bottom_in[181], chany_bottom_in[259], chany_bottom_in[277]}),
		.sram(mux_tree_tapbuf_size8_103_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_103_sram_inv[0:3]),
		.out(chanx_left_out[260]));

	mux_tree_tapbuf_size8 mux_left_track_529 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[104], chany_top_in[200], chany_bottom_in[86], chany_bottom_in[182], chany_bottom_in[263], chany_bottom_in[278]}),
		.sram(mux_tree_tapbuf_size8_104_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_104_sram_inv[0:3]),
		.out(chanx_left_out[264]));

	mux_tree_tapbuf_size8 mux_left_track_537 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[102], chany_top_in[198], chany_bottom_in[88], chany_bottom_in[184], chany_bottom_in[267], chany_bottom_in[280]}),
		.sram(mux_tree_tapbuf_size8_105_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_105_sram_inv[0:3]),
		.out(chanx_left_out[268]));

	mux_tree_tapbuf_size8 mux_left_track_545 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[101], chany_top_in[197], chany_bottom_in[89], chany_bottom_in[185], chany_bottom_in[271], chany_bottom_in[281]}),
		.sram(mux_tree_tapbuf_size8_106_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_106_sram_inv[0:3]),
		.out(chanx_left_out[272]));

	mux_tree_tapbuf_size8 mux_left_track_553 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[100], chany_top_in[196], chany_bottom_in[90], chany_bottom_in[186], chany_bottom_in[275], chany_bottom_in[282]}),
		.sram(mux_tree_tapbuf_size8_107_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_107_sram_inv[0:3]),
		.out(chanx_left_out[276]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_0_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_1_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_2_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_3_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_4_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_5_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_6_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_7_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_8_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_9_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_10_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_11_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_12_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_13_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_14_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_15_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_16_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_17_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_18_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_19_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_20_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_21_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_22_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_23_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_24_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_25_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_26_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_27_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_28_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_29_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_30_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_31_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_32_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_33_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_34_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_35_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_36_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_37_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_38_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_39_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_40_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_41_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_42_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_43_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_44_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_45_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_46_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_47_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_48_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_49_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_50_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_51_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_52_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_53_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_54_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_55_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_56_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_57_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_58_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_59_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_60_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_61_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_62_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_63_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_64_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_65_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_66_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_67_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_68_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_69_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_70_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_71_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_72_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_72_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_73_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_73_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_74_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_74_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_75_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_75_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_76_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_76_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_77_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_77_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_78_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_78_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_79_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_79_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_80_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_80_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_81_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_81_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_82_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_82_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_83_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_83_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_84_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_84_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_85_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_85_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_86_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_86_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_87_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_87_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_88_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_88_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_89_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_89_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_385 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_90_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_90_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_393 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_91_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_91_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_401 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_92_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_92_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_409 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_93_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_93_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_417 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_94_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_94_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_425 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_95_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_95_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_449 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_96_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_96_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_457 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_97_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_97_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_465 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_98_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_98_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_473 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_99_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_99_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_481 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_100_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_100_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_489 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_101_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_101_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_497 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_102_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_102_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_521 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_103_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_103_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_529 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_104_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_104_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_537 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_105_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_105_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_106_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_106_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_107_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_107_sram_inv[0:3]));

	mux_tree_tapbuf_size9 mux_bottom_track_73 (
		.in({chanx_right_in[81], chanx_right_in[177], chanx_right_in[247], chanx_right_in[273], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[13], chanx_left_in[43], chanx_left_in[109], chanx_left_in[205]}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size9 mux_bottom_track_81 (
		.in({chanx_right_in[80], chanx_right_in[176], chanx_right_in[243], chanx_right_in[272], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[14], chanx_left_in[47], chanx_left_in[110], chanx_left_in[206]}),
		.sram(mux_tree_tapbuf_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_1_sram_inv[0:3]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size9 mux_bottom_track_145 (
		.in({chanx_right_in[69], chanx_right_in[165], chanx_right_in[211], chanx_right_in[261], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[25], chanx_left_in[79], chanx_left_in[121], chanx_left_in[217]}),
		.sram(mux_tree_tapbuf_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_2_sram_inv[0:3]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size9 mux_bottom_track_153 (
		.in({chanx_right_in[68], chanx_right_in[164], chanx_right_in[207], chanx_right_in[260], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[26], chanx_left_in[83], chanx_left_in[122], chanx_left_in[218]}),
		.sram(mux_tree_tapbuf_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_3_sram_inv[0:3]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size9 mux_bottom_track_217 (
		.in({chanx_right_in[57], chanx_right_in[153], chanx_right_in[175], chanx_right_in[249], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[37], chanx_left_in[115], chanx_left_in[133], chanx_left_in[229]}),
		.sram(mux_tree_tapbuf_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_4_sram_inv[0:3]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size9 mux_bottom_track_225 (
		.in({chanx_right_in[56], chanx_right_in[152], chanx_right_in[171], chanx_right_in[248], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[38], chanx_left_in[119], chanx_left_in[134], chanx_left_in[230]}),
		.sram(mux_tree_tapbuf_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_5_sram_inv[0:3]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size9 mux_bottom_track_289 (
		.in({chanx_right_in[45], chanx_right_in[139], chanx_right_in[141], chanx_right_in[237], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[49], chanx_left_in[145], chanx_left_in[151], chanx_left_in[241]}),
		.sram(mux_tree_tapbuf_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_6_sram_inv[0:3]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size9 mux_bottom_track_297 (
		.in({chanx_right_in[44], chanx_right_in[135], chanx_right_in[140], chanx_right_in[236], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[50], chanx_left_in[146], chanx_left_in[155], chanx_left_in[242]}),
		.sram(mux_tree_tapbuf_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_7_sram_inv[0:3]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size9 mux_bottom_track_361 (
		.in({chanx_right_in[33], chanx_right_in[103], chanx_right_in[129], chanx_right_in[225], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[61], chanx_left_in[157], chanx_left_in[187], chanx_left_in[253]}),
		.sram(mux_tree_tapbuf_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_8_sram_inv[0:3]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size9 mux_bottom_track_369 (
		.in({chanx_right_in[32], chanx_right_in[99], chanx_right_in[128], chanx_right_in[224], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[62], chanx_left_in[158], chanx_left_in[191], chanx_left_in[254]}),
		.sram(mux_tree_tapbuf_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_9_sram_inv[0:3]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size9 mux_bottom_track_433 (
		.in({chanx_right_in[21], chanx_right_in[67], chanx_right_in[117], chanx_right_in[213], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[73], chanx_left_in[169], chanx_left_in[223], chanx_left_in[265]}),
		.sram(mux_tree_tapbuf_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_10_sram_inv[0:3]),
		.out(chany_bottom_out[216]));

	mux_tree_tapbuf_size9 mux_bottom_track_441 (
		.in({chanx_right_in[20], chanx_right_in[63], chanx_right_in[116], chanx_right_in[212], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[74], chanx_left_in[170], chanx_left_in[227], chanx_left_in[266]}),
		.sram(mux_tree_tapbuf_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_11_sram_inv[0:3]),
		.out(chany_bottom_out[220]));

	mux_tree_tapbuf_size9 mux_bottom_track_505 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[105], chanx_right_in[201], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[85], chanx_left_in[181], chanx_left_in[259], chanx_left_in[277]}),
		.sram(mux_tree_tapbuf_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_12_sram_inv[0:3]),
		.out(chany_bottom_out[252]));

	mux_tree_tapbuf_size9 mux_bottom_track_513 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[104], chanx_right_in[200], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[86], chanx_left_in[182], chanx_left_in[263], chanx_left_in[278]}),
		.sram(mux_tree_tapbuf_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_13_sram_inv[0:3]),
		.out(chany_bottom_out[256]));

	mux_tree_tapbuf_size9 mux_left_track_73 (
		.in({chany_top_in[84], chany_top_in[180], chany_top_in[255], chany_top_in[276], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[106], chany_bottom_in[202], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_14_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size9 mux_left_track_81 (
		.in({chany_top_in[82], chany_top_in[178], chany_top_in[251], chany_top_in[274], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[108], chany_bottom_in[204], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_15_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size9 mux_left_track_145 (
		.in({chany_top_in[72], chany_top_in[168], chany_top_in[219], chany_top_in[264], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[118], chany_bottom_in[214], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_16_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size9 mux_left_track_153 (
		.in({chany_top_in[70], chany_top_in[166], chany_top_in[215], chany_top_in[262], chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[120], chany_bottom_in[216], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_17_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size9 mux_left_track_217 (
		.in({chany_top_in[60], chany_top_in[156], chany_top_in[183], chany_top_in[252], chany_bottom_in[34], chany_bottom_in[107], chany_bottom_in[130], chany_bottom_in[226], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_18_sram_inv[0:3]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size9 mux_left_track_225 (
		.in({chany_top_in[58], chany_top_in[154], chany_top_in[179], chany_top_in[250], chany_bottom_in[36], chany_bottom_in[111], chany_bottom_in[132], chany_bottom_in[228], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_19_sram_inv[0:3]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size9 mux_left_track_289 (
		.in({chany_top_in[48], chany_top_in[144], chany_top_in[147], chany_top_in[240], chany_bottom_in[46], chany_bottom_in[142:143], chany_bottom_in[238], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_20_sram_inv[0:3]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size9 mux_left_track_297 (
		.in({chany_top_in[46], chany_top_in[142:143], chany_top_in[238], chany_bottom_in[48], chany_bottom_in[144], chany_bottom_in[147], chany_bottom_in[240], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_21_sram_inv[0:3]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size9 mux_left_track_361 (
		.in({chany_top_in[36], chany_top_in[111], chany_top_in[132], chany_top_in[228], chany_bottom_in[58], chany_bottom_in[154], chany_bottom_in[179], chany_bottom_in[250], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_22_sram_inv[0:3]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size9 mux_left_track_369 (
		.in({chany_top_in[34], chany_top_in[107], chany_top_in[130], chany_top_in[226], chany_bottom_in[60], chany_bottom_in[156], chany_bottom_in[183], chany_bottom_in[252], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_23_sram_inv[0:3]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size9 mux_left_track_433 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[120], chany_top_in[216], chany_bottom_in[70], chany_bottom_in[166], chany_bottom_in[215], chany_bottom_in[262], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_24_sram_inv[0:3]),
		.out(chanx_left_out[216]));

	mux_tree_tapbuf_size9 mux_left_track_441 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[118], chany_top_in[214], chany_bottom_in[72], chany_bottom_in[168], chany_bottom_in[219], chany_bottom_in[264], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_25_sram_inv[0:3]),
		.out(chanx_left_out[220]));

	mux_tree_tapbuf_size9 mux_left_track_505 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[108], chany_top_in[204], chany_bottom_in[82], chany_bottom_in[178], chany_bottom_in[251], chany_bottom_in[274], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_26_sram_inv[0:3]),
		.out(chanx_left_out[252]));

	mux_tree_tapbuf_size9 mux_left_track_513 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[106], chany_top_in[202], chany_bottom_in[84], chany_bottom_in[180], chany_bottom_in[255], chany_bottom_in[276], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_27_sram_inv[0:3]),
		.out(chanx_left_out[256]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_18_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_19_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_20_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_21_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_22_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_23_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_433 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_24_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_441 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_25_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_505 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_26_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_513 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_27_sram_inv[0:3]));

	mux_tree_tapbuf_size7 mux_bottom_track_545 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[98], chanx_right_in[194], chanx_left_in[92], chanx_left_in[188], chanx_left_in[279]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[272]));

	mux_tree_tapbuf_size7 mux_bottom_track_553 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[97], chanx_right_in[193], chanx_left_in[93], chanx_left_in[189], chanx_left_in[283]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[276]));

	mux_tree_tapbuf_size7 mux_bottom_track_561 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[96], chanx_right_in[192], chanx_left_in[94], chanx_left_in[190], chanx_left_in[284]}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[280]));

	mux_tree_tapbuf_size7 mux_bottom_track_569 (
		.in({chanx_right_in[94], chanx_right_in[190], chanx_right_in[284], chanx_left_in[0], chanx_left_in[3], chanx_left_in[96], chanx_left_in[192]}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[284]));

	mux_tree_tapbuf_size7 mux_left_track_17 (
		.in({chany_top_in[93], chany_top_in[189], chany_top_in[283], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[97], chany_bottom_in[193]}),
		.sram(mux_tree_tapbuf_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_4_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size7 mux_left_track_25 (
		.in({chany_top_in[92], chany_top_in[188], chany_top_in[279], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[98], chany_bottom_in[194]}),
		.sram(mux_tree_tapbuf_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_5_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size7 mux_left_track_561 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[98], chany_top_in[194], chany_bottom_in[92], chany_bottom_in[188], chany_bottom_in[279]}),
		.sram(mux_tree_tapbuf_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_6_sram_inv[0:2]),
		.out(chanx_left_out[280]));

	mux_tree_tapbuf_size7 mux_left_track_569 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[97], chany_top_in[193], chany_bottom_in[93], chany_bottom_in[189], chany_bottom_in[283]}),
		.sram(mux_tree_tapbuf_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_7_sram_inv[0:2]),
		.out(chanx_left_out[284]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_545 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_553 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_561 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_569 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_7_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_5__5_ -----

//----- Default net type -----
`default_nettype wire



