//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[4][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Jun 27 10:27:38 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_4__2_ -----
module sb_4__2_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_,
                ccff_head,
                chany_top_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:188] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:188] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
//----- INPUT PORTS -----
input [0:188] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:188] chany_top_out;
//----- OUTPUT PORTS -----
output [0:188] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:188] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_1_sram;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_2_sram;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_3_sram;
wire [0:3] mux_tree_tapbuf_size10_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_3_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_11_sram;
wire [0:3] mux_tree_tapbuf_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_12_sram;
wire [0:3] mux_tree_tapbuf_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_13_sram;
wire [0:3] mux_tree_tapbuf_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_14_sram;
wire [0:3] mux_tree_tapbuf_size11_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_15_sram;
wire [0:3] mux_tree_tapbuf_size11_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_16_sram;
wire [0:3] mux_tree_tapbuf_size11_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_17_sram;
wire [0:3] mux_tree_tapbuf_size11_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_18_sram;
wire [0:3] mux_tree_tapbuf_size11_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_19_sram;
wire [0:3] mux_tree_tapbuf_size11_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_20_sram;
wire [0:3] mux_tree_tapbuf_size11_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_21_sram;
wire [0:3] mux_tree_tapbuf_size11_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_22_sram;
wire [0:3] mux_tree_tapbuf_size11_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_23_sram;
wire [0:3] mux_tree_tapbuf_size11_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_24_sram;
wire [0:3] mux_tree_tapbuf_size11_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_25_sram;
wire [0:3] mux_tree_tapbuf_size11_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_26_sram;
wire [0:3] mux_tree_tapbuf_size11_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_27_sram;
wire [0:3] mux_tree_tapbuf_size11_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_28_sram;
wire [0:3] mux_tree_tapbuf_size11_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_29_sram;
wire [0:3] mux_tree_tapbuf_size11_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_30_sram;
wire [0:3] mux_tree_tapbuf_size11_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_31_sram;
wire [0:3] mux_tree_tapbuf_size11_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_32_sram;
wire [0:3] mux_tree_tapbuf_size11_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_33_sram;
wire [0:3] mux_tree_tapbuf_size11_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_34_sram;
wire [0:3] mux_tree_tapbuf_size11_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_35_sram;
wire [0:3] mux_tree_tapbuf_size11_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_36_sram;
wire [0:3] mux_tree_tapbuf_size11_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_37_sram;
wire [0:3] mux_tree_tapbuf_size11_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_38_sram;
wire [0:3] mux_tree_tapbuf_size11_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_39_sram;
wire [0:3] mux_tree_tapbuf_size11_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_40_sram;
wire [0:3] mux_tree_tapbuf_size11_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_41_sram;
wire [0:3] mux_tree_tapbuf_size11_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_42_sram;
wire [0:3] mux_tree_tapbuf_size11_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_43_sram;
wire [0:3] mux_tree_tapbuf_size11_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_44_sram;
wire [0:3] mux_tree_tapbuf_size11_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_45_sram;
wire [0:3] mux_tree_tapbuf_size11_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_46_sram;
wire [0:3] mux_tree_tapbuf_size11_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_47_sram;
wire [0:3] mux_tree_tapbuf_size11_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_48_sram;
wire [0:3] mux_tree_tapbuf_size11_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_49_sram;
wire [0:3] mux_tree_tapbuf_size11_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_50_sram;
wire [0:3] mux_tree_tapbuf_size11_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_51_sram;
wire [0:3] mux_tree_tapbuf_size11_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_100_sram;
wire [0:3] mux_tree_tapbuf_size12_100_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_101_sram;
wire [0:3] mux_tree_tapbuf_size12_101_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_102_sram;
wire [0:3] mux_tree_tapbuf_size12_102_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_103_sram;
wire [0:3] mux_tree_tapbuf_size12_103_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_104_sram;
wire [0:3] mux_tree_tapbuf_size12_104_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_105_sram;
wire [0:3] mux_tree_tapbuf_size12_105_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_106_sram;
wire [0:3] mux_tree_tapbuf_size12_106_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_107_sram;
wire [0:3] mux_tree_tapbuf_size12_107_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_108_sram;
wire [0:3] mux_tree_tapbuf_size12_108_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_109_sram;
wire [0:3] mux_tree_tapbuf_size12_109_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_110_sram;
wire [0:3] mux_tree_tapbuf_size12_110_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_111_sram;
wire [0:3] mux_tree_tapbuf_size12_111_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_112_sram;
wire [0:3] mux_tree_tapbuf_size12_112_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_113_sram;
wire [0:3] mux_tree_tapbuf_size12_113_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_114_sram;
wire [0:3] mux_tree_tapbuf_size12_114_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_115_sram;
wire [0:3] mux_tree_tapbuf_size12_115_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_116_sram;
wire [0:3] mux_tree_tapbuf_size12_116_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_117_sram;
wire [0:3] mux_tree_tapbuf_size12_117_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_118_sram;
wire [0:3] mux_tree_tapbuf_size12_118_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_119_sram;
wire [0:3] mux_tree_tapbuf_size12_119_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_120_sram;
wire [0:3] mux_tree_tapbuf_size12_120_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_121_sram;
wire [0:3] mux_tree_tapbuf_size12_121_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_122_sram;
wire [0:3] mux_tree_tapbuf_size12_122_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_123_sram;
wire [0:3] mux_tree_tapbuf_size12_123_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_124_sram;
wire [0:3] mux_tree_tapbuf_size12_124_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_125_sram;
wire [0:3] mux_tree_tapbuf_size12_125_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_126_sram;
wire [0:3] mux_tree_tapbuf_size12_126_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_127_sram;
wire [0:3] mux_tree_tapbuf_size12_127_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_128_sram;
wire [0:3] mux_tree_tapbuf_size12_128_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_129_sram;
wire [0:3] mux_tree_tapbuf_size12_129_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_130_sram;
wire [0:3] mux_tree_tapbuf_size12_130_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_131_sram;
wire [0:3] mux_tree_tapbuf_size12_131_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_132_sram;
wire [0:3] mux_tree_tapbuf_size12_132_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_36_sram;
wire [0:3] mux_tree_tapbuf_size12_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_37_sram;
wire [0:3] mux_tree_tapbuf_size12_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_38_sram;
wire [0:3] mux_tree_tapbuf_size12_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_39_sram;
wire [0:3] mux_tree_tapbuf_size12_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_40_sram;
wire [0:3] mux_tree_tapbuf_size12_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_41_sram;
wire [0:3] mux_tree_tapbuf_size12_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_42_sram;
wire [0:3] mux_tree_tapbuf_size12_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_43_sram;
wire [0:3] mux_tree_tapbuf_size12_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_44_sram;
wire [0:3] mux_tree_tapbuf_size12_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_45_sram;
wire [0:3] mux_tree_tapbuf_size12_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_46_sram;
wire [0:3] mux_tree_tapbuf_size12_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_47_sram;
wire [0:3] mux_tree_tapbuf_size12_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_48_sram;
wire [0:3] mux_tree_tapbuf_size12_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_49_sram;
wire [0:3] mux_tree_tapbuf_size12_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_50_sram;
wire [0:3] mux_tree_tapbuf_size12_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_51_sram;
wire [0:3] mux_tree_tapbuf_size12_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_52_sram;
wire [0:3] mux_tree_tapbuf_size12_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_53_sram;
wire [0:3] mux_tree_tapbuf_size12_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_54_sram;
wire [0:3] mux_tree_tapbuf_size12_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_55_sram;
wire [0:3] mux_tree_tapbuf_size12_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_56_sram;
wire [0:3] mux_tree_tapbuf_size12_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_57_sram;
wire [0:3] mux_tree_tapbuf_size12_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_58_sram;
wire [0:3] mux_tree_tapbuf_size12_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_59_sram;
wire [0:3] mux_tree_tapbuf_size12_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_60_sram;
wire [0:3] mux_tree_tapbuf_size12_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_61_sram;
wire [0:3] mux_tree_tapbuf_size12_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_62_sram;
wire [0:3] mux_tree_tapbuf_size12_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_63_sram;
wire [0:3] mux_tree_tapbuf_size12_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_64_sram;
wire [0:3] mux_tree_tapbuf_size12_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_65_sram;
wire [0:3] mux_tree_tapbuf_size12_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_66_sram;
wire [0:3] mux_tree_tapbuf_size12_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_67_sram;
wire [0:3] mux_tree_tapbuf_size12_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_68_sram;
wire [0:3] mux_tree_tapbuf_size12_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_69_sram;
wire [0:3] mux_tree_tapbuf_size12_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_70_sram;
wire [0:3] mux_tree_tapbuf_size12_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_71_sram;
wire [0:3] mux_tree_tapbuf_size12_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_72_sram;
wire [0:3] mux_tree_tapbuf_size12_72_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_73_sram;
wire [0:3] mux_tree_tapbuf_size12_73_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_74_sram;
wire [0:3] mux_tree_tapbuf_size12_74_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_75_sram;
wire [0:3] mux_tree_tapbuf_size12_75_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_76_sram;
wire [0:3] mux_tree_tapbuf_size12_76_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_77_sram;
wire [0:3] mux_tree_tapbuf_size12_77_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_78_sram;
wire [0:3] mux_tree_tapbuf_size12_78_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_79_sram;
wire [0:3] mux_tree_tapbuf_size12_79_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_80_sram;
wire [0:3] mux_tree_tapbuf_size12_80_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_81_sram;
wire [0:3] mux_tree_tapbuf_size12_81_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_82_sram;
wire [0:3] mux_tree_tapbuf_size12_82_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_83_sram;
wire [0:3] mux_tree_tapbuf_size12_83_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_84_sram;
wire [0:3] mux_tree_tapbuf_size12_84_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_85_sram;
wire [0:3] mux_tree_tapbuf_size12_85_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_86_sram;
wire [0:3] mux_tree_tapbuf_size12_86_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_87_sram;
wire [0:3] mux_tree_tapbuf_size12_87_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_88_sram;
wire [0:3] mux_tree_tapbuf_size12_88_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_89_sram;
wire [0:3] mux_tree_tapbuf_size12_89_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_90_sram;
wire [0:3] mux_tree_tapbuf_size12_90_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_91_sram;
wire [0:3] mux_tree_tapbuf_size12_91_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_92_sram;
wire [0:3] mux_tree_tapbuf_size12_92_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_93_sram;
wire [0:3] mux_tree_tapbuf_size12_93_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_94_sram;
wire [0:3] mux_tree_tapbuf_size12_94_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_95_sram;
wire [0:3] mux_tree_tapbuf_size12_95_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_96_sram;
wire [0:3] mux_tree_tapbuf_size12_96_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_97_sram;
wire [0:3] mux_tree_tapbuf_size12_97_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_98_sram;
wire [0:3] mux_tree_tapbuf_size12_98_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_99_sram;
wire [0:3] mux_tree_tapbuf_size12_99_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size15_0_sram;
wire [0:3] mux_tree_tapbuf_size15_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_1_sram;
wire [0:3] mux_tree_tapbuf_size15_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_2_sram;
wire [0:3] mux_tree_tapbuf_size15_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_2_ccff_tail;
wire [0:4] mux_tree_tapbuf_size16_0_sram;
wire [0:4] mux_tree_tapbuf_size16_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_10_sram;
wire [0:4] mux_tree_tapbuf_size16_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_11_sram;
wire [0:4] mux_tree_tapbuf_size16_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_12_sram;
wire [0:4] mux_tree_tapbuf_size16_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_13_sram;
wire [0:4] mux_tree_tapbuf_size16_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_14_sram;
wire [0:4] mux_tree_tapbuf_size16_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_15_sram;
wire [0:4] mux_tree_tapbuf_size16_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_16_sram;
wire [0:4] mux_tree_tapbuf_size16_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_17_sram;
wire [0:4] mux_tree_tapbuf_size16_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_18_sram;
wire [0:4] mux_tree_tapbuf_size16_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_19_sram;
wire [0:4] mux_tree_tapbuf_size16_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_1_sram;
wire [0:4] mux_tree_tapbuf_size16_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_20_sram;
wire [0:4] mux_tree_tapbuf_size16_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_21_sram;
wire [0:4] mux_tree_tapbuf_size16_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_22_sram;
wire [0:4] mux_tree_tapbuf_size16_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_23_sram;
wire [0:4] mux_tree_tapbuf_size16_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_24_sram;
wire [0:4] mux_tree_tapbuf_size16_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_25_sram;
wire [0:4] mux_tree_tapbuf_size16_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_26_sram;
wire [0:4] mux_tree_tapbuf_size16_26_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_27_sram;
wire [0:4] mux_tree_tapbuf_size16_27_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_28_sram;
wire [0:4] mux_tree_tapbuf_size16_28_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_29_sram;
wire [0:4] mux_tree_tapbuf_size16_29_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_2_sram;
wire [0:4] mux_tree_tapbuf_size16_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_30_sram;
wire [0:4] mux_tree_tapbuf_size16_30_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_31_sram;
wire [0:4] mux_tree_tapbuf_size16_31_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_32_sram;
wire [0:4] mux_tree_tapbuf_size16_32_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_33_sram;
wire [0:4] mux_tree_tapbuf_size16_33_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_34_sram;
wire [0:4] mux_tree_tapbuf_size16_34_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_35_sram;
wire [0:4] mux_tree_tapbuf_size16_35_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_36_sram;
wire [0:4] mux_tree_tapbuf_size16_36_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_37_sram;
wire [0:4] mux_tree_tapbuf_size16_37_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_38_sram;
wire [0:4] mux_tree_tapbuf_size16_38_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_39_sram;
wire [0:4] mux_tree_tapbuf_size16_39_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_3_sram;
wire [0:4] mux_tree_tapbuf_size16_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_40_sram;
wire [0:4] mux_tree_tapbuf_size16_40_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_41_sram;
wire [0:4] mux_tree_tapbuf_size16_41_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_42_sram;
wire [0:4] mux_tree_tapbuf_size16_42_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_43_sram;
wire [0:4] mux_tree_tapbuf_size16_43_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_44_sram;
wire [0:4] mux_tree_tapbuf_size16_44_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_4_sram;
wire [0:4] mux_tree_tapbuf_size16_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_5_sram;
wire [0:4] mux_tree_tapbuf_size16_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_6_sram;
wire [0:4] mux_tree_tapbuf_size16_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_7_sram;
wire [0:4] mux_tree_tapbuf_size16_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_8_sram;
wire [0:4] mux_tree_tapbuf_size16_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size16_9_sram;
wire [0:4] mux_tree_tapbuf_size16_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size16_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size16_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_25_sram;
wire [0:2] mux_tree_tapbuf_size5_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_26_sram;
wire [0:2] mux_tree_tapbuf_size5_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_27_sram;
wire [0:2] mux_tree_tapbuf_size5_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_28_sram;
wire [0:2] mux_tree_tapbuf_size5_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_29_sram;
wire [0:2] mux_tree_tapbuf_size5_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_30_sram;
wire [0:2] mux_tree_tapbuf_size5_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_31_sram;
wire [0:2] mux_tree_tapbuf_size5_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_32_sram;
wire [0:2] mux_tree_tapbuf_size5_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_33_sram;
wire [0:2] mux_tree_tapbuf_size5_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_34_sram;
wire [0:2] mux_tree_tapbuf_size5_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_35_sram;
wire [0:2] mux_tree_tapbuf_size5_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_36_sram;
wire [0:2] mux_tree_tapbuf_size5_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_37_sram;
wire [0:2] mux_tree_tapbuf_size5_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_38_sram;
wire [0:2] mux_tree_tapbuf_size5_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_39_sram;
wire [0:2] mux_tree_tapbuf_size5_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_40_sram;
wire [0:2] mux_tree_tapbuf_size5_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_41_sram;
wire [0:2] mux_tree_tapbuf_size5_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_42_sram;
wire [0:2] mux_tree_tapbuf_size5_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_43_sram;
wire [0:2] mux_tree_tapbuf_size5_43_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_44_sram;
wire [0:2] mux_tree_tapbuf_size5_44_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size6 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[0], chanx_left_in[48], chanx_left_in[96], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size6 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[44], chanx_left_in[92], chanx_left_in[140], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size6 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[43], chanx_left_in[91], chanx_left_in[139], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size6_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[47], chanx_left_in[95], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size5 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[46], chanx_left_in[94], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size5 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[45], chanx_left_in[93], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size5 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[42], chanx_left_in[90], chanx_left_in[138], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size5 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[41], chanx_left_in[89], chanx_left_in[137], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size5 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[40], chanx_left_in[88], chanx_left_in[136], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size5 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[39], chanx_left_in[87], chanx_left_in[135], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size5 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[38], chanx_left_in[86], chanx_left_in[134], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size5 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[37], chanx_left_in[85], chanx_left_in[133], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size5 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[36], chanx_left_in[84], chanx_left_in[132], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size5 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[35], chanx_left_in[83], chanx_left_in[131], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size5 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[34], chanx_left_in[82], chanx_left_in[130], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size5 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[33], chanx_left_in[81], chanx_left_in[129], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size5 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[32], chanx_left_in[80], chanx_left_in[128], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size5 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[31], chanx_left_in[79], chanx_left_in[127], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size5 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[30], chanx_left_in[78], chanx_left_in[126], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size5 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[29], chanx_left_in[77], chanx_left_in[125], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size5 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[28], chanx_left_in[76], chanx_left_in[124], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size5 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[27], chanx_left_in[75], chanx_left_in[123], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size5 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[26], chanx_left_in[74], chanx_left_in[122], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size5 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[25], chanx_left_in[73], chanx_left_in[121], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size5 mux_top_track_192 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[24], chanx_left_in[72], chanx_left_in[120], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size5 mux_top_track_200 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[23], chanx_left_in[71], chanx_left_in[119], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size5 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[22], chanx_left_in[70], chanx_left_in[118], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size5 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[21], chanx_left_in[69], chanx_left_in[117], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size5 mux_top_track_224 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[20], chanx_left_in[68], chanx_left_in[116], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size5_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_25_sram_inv[0:2]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size5 mux_top_track_232 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[19], chanx_left_in[67], chanx_left_in[115], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size5_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_26_sram_inv[0:2]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size5 mux_top_track_240 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[18], chanx_left_in[66], chanx_left_in[114], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size5_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_27_sram_inv[0:2]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size5 mux_top_track_248 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[17], chanx_left_in[65], chanx_left_in[113], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size5_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_28_sram_inv[0:2]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size5 mux_top_track_256 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[16], chanx_left_in[64], chanx_left_in[112], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size5_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_29_sram_inv[0:2]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size5 mux_top_track_264 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[15], chanx_left_in[63], chanx_left_in[111], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size5_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_30_sram_inv[0:2]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size5 mux_top_track_272 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[14], chanx_left_in[62], chanx_left_in[110], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size5_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_31_sram_inv[0:2]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size5 mux_top_track_280 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[13], chanx_left_in[61], chanx_left_in[109], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size5_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_32_sram_inv[0:2]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size5 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[12], chanx_left_in[60], chanx_left_in[108], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size5_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_33_sram_inv[0:2]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size5 mux_top_track_296 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[11], chanx_left_in[59], chanx_left_in[107], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size5_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_34_sram_inv[0:2]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size5 mux_top_track_304 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[10], chanx_left_in[58], chanx_left_in[106], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size5_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_35_sram_inv[0:2]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size5 mux_top_track_312 (
		.in({top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[9], chanx_left_in[57], chanx_left_in[105], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size5_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_36_sram_inv[0:2]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size5 mux_top_track_320 (
		.in({top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[8], chanx_left_in[56], chanx_left_in[104], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size5_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_37_sram_inv[0:2]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size5 mux_top_track_328 (
		.in({top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[7], chanx_left_in[55], chanx_left_in[103], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size5_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_38_sram_inv[0:2]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size5 mux_top_track_336 (
		.in({top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[6], chanx_left_in[54], chanx_left_in[102], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size5_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_39_sram_inv[0:2]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size5 mux_top_track_344 (
		.in({top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[5], chanx_left_in[53], chanx_left_in[101], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size5_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_40_sram_inv[0:2]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size5 mux_top_track_352 (
		.in({top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[4], chanx_left_in[52], chanx_left_in[100], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size5_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_41_sram_inv[0:2]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size5 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[3], chanx_left_in[51], chanx_left_in[99], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size5_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_42_sram_inv[0:2]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size5 mux_top_track_368 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[2], chanx_left_in[50], chanx_left_in[98], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size5_43_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_43_sram_inv[0:2]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size5 mux_top_track_376 (
		.in({top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[1], chanx_left_in[49], chanx_left_in[97], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size5_44_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_44_sram_inv[0:2]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size5_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_25_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_26_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_27_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_28_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_29_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_30_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_31_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_32_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_33_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_34_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_35_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_36_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_37_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_38_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_39_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_40_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_41_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_42_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_43_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_43_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_44_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_44_sram_inv[0:2]));

	mux_tree_tapbuf_size16 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[1], chanx_left_in[49], chanx_left_in[97], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size16_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_0_sram_inv[0:4]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size16 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[2], chanx_left_in[50], chanx_left_in[98], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size16_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_1_sram_inv[0:4]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size16 mux_bottom_track_17 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[3], chanx_left_in[51], chanx_left_in[99], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size16_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_2_sram_inv[0:4]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size16 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[4], chanx_left_in[52], chanx_left_in[100], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size16_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_3_sram_inv[0:4]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size16 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[5], chanx_left_in[53], chanx_left_in[101], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size16_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_4_sram_inv[0:4]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size16 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[6], chanx_left_in[54], chanx_left_in[102], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size16_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_5_sram_inv[0:4]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size16 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[7], chanx_left_in[55], chanx_left_in[103], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size16_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_6_sram_inv[0:4]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size16 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[8], chanx_left_in[56], chanx_left_in[104], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size16_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_7_sram_inv[0:4]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size16 mux_bottom_track_65 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[9], chanx_left_in[57], chanx_left_in[105], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size16_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_8_sram_inv[0:4]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size16 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[10], chanx_left_in[58], chanx_left_in[106], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size16_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_9_sram_inv[0:4]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size16 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[11], chanx_left_in[59], chanx_left_in[107], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size16_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_10_sram_inv[0:4]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size16 mux_bottom_track_89 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[12], chanx_left_in[60], chanx_left_in[108], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size16_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_11_sram_inv[0:4]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size16 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[13], chanx_left_in[61], chanx_left_in[109], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size16_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_12_sram_inv[0:4]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size16 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[14], chanx_left_in[62], chanx_left_in[110], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size16_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_13_sram_inv[0:4]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size16 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[15], chanx_left_in[63], chanx_left_in[111], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size16_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_14_sram_inv[0:4]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size16 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[16], chanx_left_in[64], chanx_left_in[112], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size16_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_15_sram_inv[0:4]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size16 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[17], chanx_left_in[65], chanx_left_in[113], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size16_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_16_sram_inv[0:4]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size16 mux_bottom_track_137 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[18], chanx_left_in[66], chanx_left_in[114], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size16_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_17_sram_inv[0:4]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size16 mux_bottom_track_145 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[19], chanx_left_in[67], chanx_left_in[115], chanx_left_in[163]}),
		.sram(mux_tree_tapbuf_size16_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_18_sram_inv[0:4]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size16 mux_bottom_track_153 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[20], chanx_left_in[68], chanx_left_in[116], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size16_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_19_sram_inv[0:4]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size16 mux_bottom_track_161 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[21], chanx_left_in[69], chanx_left_in[117], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size16_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_20_sram_inv[0:4]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size16 mux_bottom_track_169 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[22], chanx_left_in[70], chanx_left_in[118], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size16_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_21_sram_inv[0:4]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size16 mux_bottom_track_177 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[23], chanx_left_in[71], chanx_left_in[119], chanx_left_in[167]}),
		.sram(mux_tree_tapbuf_size16_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_22_sram_inv[0:4]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size16 mux_bottom_track_185 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[24], chanx_left_in[72], chanx_left_in[120], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size16_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_23_sram_inv[0:4]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size16 mux_bottom_track_193 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[25], chanx_left_in[73], chanx_left_in[121], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size16_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_24_sram_inv[0:4]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size16 mux_bottom_track_201 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[26], chanx_left_in[74], chanx_left_in[122], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size16_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_25_sram_inv[0:4]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size16 mux_bottom_track_209 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[27], chanx_left_in[75], chanx_left_in[123], chanx_left_in[171]}),
		.sram(mux_tree_tapbuf_size16_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_26_sram_inv[0:4]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size16 mux_bottom_track_217 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[28], chanx_left_in[76], chanx_left_in[124], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size16_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_27_sram_inv[0:4]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size16 mux_bottom_track_225 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[29], chanx_left_in[77], chanx_left_in[125], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size16_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_28_sram_inv[0:4]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size16 mux_bottom_track_233 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[30], chanx_left_in[78], chanx_left_in[126], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size16_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_29_sram_inv[0:4]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size16 mux_bottom_track_241 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[31], chanx_left_in[79], chanx_left_in[127], chanx_left_in[175]}),
		.sram(mux_tree_tapbuf_size16_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_30_sram_inv[0:4]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size16 mux_bottom_track_249 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[32], chanx_left_in[80], chanx_left_in[128], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size16_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_31_sram_inv[0:4]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size16 mux_bottom_track_257 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[33], chanx_left_in[81], chanx_left_in[129], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size16_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_32_sram_inv[0:4]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size16 mux_bottom_track_265 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[34], chanx_left_in[82], chanx_left_in[130], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size16_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_33_sram_inv[0:4]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size16 mux_bottom_track_273 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[35], chanx_left_in[83], chanx_left_in[131], chanx_left_in[179]}),
		.sram(mux_tree_tapbuf_size16_34_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_34_sram_inv[0:4]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size16 mux_bottom_track_281 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[36], chanx_left_in[84], chanx_left_in[132], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size16_35_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_35_sram_inv[0:4]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size16 mux_bottom_track_289 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[37], chanx_left_in[85], chanx_left_in[133], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size16_36_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_36_sram_inv[0:4]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size16 mux_bottom_track_297 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[38], chanx_left_in[86], chanx_left_in[134], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size16_37_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_37_sram_inv[0:4]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size16 mux_bottom_track_305 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[39], chanx_left_in[87], chanx_left_in[135], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size16_38_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_38_sram_inv[0:4]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size16 mux_bottom_track_313 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[40], chanx_left_in[88], chanx_left_in[136], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size16_39_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_39_sram_inv[0:4]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size16 mux_bottom_track_321 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[41], chanx_left_in[89], chanx_left_in[137], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size16_40_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_40_sram_inv[0:4]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size16 mux_bottom_track_329 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[42], chanx_left_in[90], chanx_left_in[138], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size16_41_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_41_sram_inv[0:4]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size16 mux_bottom_track_337 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[43], chanx_left_in[91], chanx_left_in[139], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size16_42_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_42_sram_inv[0:4]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size16 mux_bottom_track_345 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[44], chanx_left_in[92], chanx_left_in[140], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size16_43_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_43_sram_inv[0:4]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size16 mux_bottom_track_377 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[0], chanx_left_in[48], chanx_left_in[96], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size16_44_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size16_44_sram_inv[0:4]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_0_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_1_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_2_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_3_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_4_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_5_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_6_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_7_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_8_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_9_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_10_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_11_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_12_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_13_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_14_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_15_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_16_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_17_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_18_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_19_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_20_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_21_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_22_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_23_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_24_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_25_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_26_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_27_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_28_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_29_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_30_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_31_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_32_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_33_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_34_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_34_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_35_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_35_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_36_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_36_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_37_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_37_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_38_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_38_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_39_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_39_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_40_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_40_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_41_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_41_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_42_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_42_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_43_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_43_sram_inv[0:4]));

	mux_tree_tapbuf_size16_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size16_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size16_44_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size16_44_sram_inv[0:4]));

	mux_tree_tapbuf_size15 mux_bottom_track_353 (
		.in({bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[45], chanx_left_in[93], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size15_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_0_sram_inv[0:3]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size15 mux_bottom_track_361 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[46], chanx_left_in[94], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size15_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_1_sram_inv[0:3]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size15 mux_bottom_track_369 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[47], chanx_left_in[95], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size15_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_2_sram_inv[0:3]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size15_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_0_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_1_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size12 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[3], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size12 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[7], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size12 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size12 mux_left_track_9 (
		.in({chany_bottom_in[4], chany_bottom_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size12 mux_left_track_11 (
		.in({chany_bottom_in[5], chany_bottom_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size12 mux_left_track_13 (
		.in({chany_bottom_in[6], chany_bottom_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size12 mux_left_track_19 (
		.in({chany_bottom_in[10], chany_bottom_in[35], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size12 mux_left_track_21 (
		.in({chany_bottom_in[12], chany_bottom_in[39], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size12 mux_left_track_23 (
		.in({chany_bottom_in[13], chany_bottom_in[43], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size12 mux_left_track_25 (
		.in({chany_bottom_in[14], chany_bottom_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size12 mux_left_track_27 (
		.in({chany_bottom_in[16], chany_bottom_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size12 mux_left_track_29 (
		.in({chany_bottom_in[17], chany_bottom_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size12 mux_left_track_31 (
		.in({chany_bottom_in[18], chany_bottom_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size12 mux_left_track_37 (
		.in({chany_bottom_in[22], chany_bottom_in[71], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size12 mux_left_track_39 (
		.in({chany_bottom_in[24], chany_bottom_in[75], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size12 mux_left_track_41 (
		.in({chany_bottom_in[25], chany_bottom_in[79], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size12 mux_left_track_43 (
		.in({chany_bottom_in[26], chany_bottom_in[83], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size12 mux_left_track_45 (
		.in({chany_bottom_in[28], chany_bottom_in[87], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size12 mux_left_track_47 (
		.in({chany_bottom_in[29], chany_bottom_in[91], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size12 mux_left_track_49 (
		.in({chany_bottom_in[30], chany_bottom_in[95], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size12 mux_left_track_57 (
		.in({chany_bottom_in[36], chany_bottom_in[111], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size12 mux_left_track_59 (
		.in({chany_bottom_in[37], chany_bottom_in[115], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size12 mux_left_track_61 (
		.in({chany_bottom_in[38], chany_bottom_in[119], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size12 mux_left_track_63 (
		.in({chany_bottom_in[40], chany_bottom_in[123], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size12 mux_left_track_65 (
		.in({chany_bottom_in[41], chany_bottom_in[127], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size12 mux_left_track_67 (
		.in({chany_bottom_in[42], chany_bottom_in[131], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size12 mux_left_track_73 (
		.in({chany_bottom_in[46], chany_bottom_in[143], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size12 mux_left_track_77 (
		.in({chany_bottom_in[49], chany_bottom_in[151], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size12 mux_left_track_79 (
		.in({chany_bottom_in[50], chany_bottom_in[155], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size12 mux_left_track_81 (
		.in({chany_bottom_in[52], chany_bottom_in[159], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size12 mux_left_track_83 (
		.in({chany_bottom_in[53], chany_bottom_in[163], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size12 mux_left_track_85 (
		.in({chany_bottom_in[54], chany_bottom_in[167], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size12 mux_left_track_91 (
		.in({chany_bottom_in[58], chany_bottom_in[179], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size12 mux_left_track_93 (
		.in({chany_bottom_in[60], chany_bottom_in[183], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size12 mux_left_track_97 (
		.in({chany_bottom_in[62], chany_bottom_in[188], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size12 mux_left_track_99 (
		.in({chany_top_in[186], chany_bottom_in[64], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_36_sram_inv[0:3]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size12 mux_left_track_101 (
		.in({chany_top_in[185], chany_bottom_in[65], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_37_sram_inv[0:3]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size12 mux_left_track_103 (
		.in({chany_top_in[184], chany_bottom_in[66], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_38_sram_inv[0:3]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size12 mux_left_track_109 (
		.in({chany_top_in[180], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_39_sram_inv[0:3]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size12 mux_left_track_111 (
		.in({chany_top_in[178], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_40_sram_inv[0:3]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size12 mux_left_track_113 (
		.in({chany_top_in[177], chany_bottom_in[73], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_41_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size12 mux_left_track_117 (
		.in({chany_top_in[174], chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_42_sram_inv[0:3]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size12 mux_left_track_119 (
		.in({chany_top_in[173], chany_bottom_in[77], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_43_sram_inv[0:3]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size12 mux_left_track_121 (
		.in({chany_top_in[172], chany_bottom_in[78], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_44_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size12 mux_left_track_127 (
		.in({chany_top_in[168], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_45_sram_inv[0:3]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size12 mux_left_track_129 (
		.in({chany_top_in[166], chany_bottom_in[84], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_46_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size12 mux_left_track_131 (
		.in({chany_top_in[165], chany_bottom_in[85], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_47_sram_inv[0:3]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size12 mux_left_track_133 (
		.in({chany_top_in[164], chany_bottom_in[86], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_48_sram_inv[0:3]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size12 mux_left_track_137 (
		.in({chany_top_in[161], chany_bottom_in[89], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_49_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size12 mux_left_track_139 (
		.in({chany_top_in[160], chany_bottom_in[90], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_50_sram_inv[0:3]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size12 mux_left_track_145 (
		.in({chany_top_in[156], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_51_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size12 mux_left_track_147 (
		.in({chany_top_in[154], chany_bottom_in[96], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_52_sram_inv[0:3]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_size12 mux_left_track_149 (
		.in({chany_top_in[153], chany_bottom_in[97], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_53_sram_inv[0:3]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_size12 mux_left_track_151 (
		.in({chany_top_in[152], chany_bottom_in[98], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_54_sram_inv[0:3]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_size12 mux_left_track_153 (
		.in({chany_top_in[150], chany_bottom_in[100], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_55_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size12 mux_left_track_155 (
		.in({chany_top_in[149], chany_bottom_in[101], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_56_sram_inv[0:3]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_size12 mux_left_track_157 (
		.in({chany_top_in[148], chany_bottom_in[102], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_57_sram_inv[0:3]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_size12 mux_left_track_163 (
		.in({chany_top_in[144], chany_bottom_in[106], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_58_sram_inv[0:3]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_size12 mux_left_track_165 (
		.in({chany_top_in[142], chany_bottom_in[108], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_59_sram_inv[0:3]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_size12 mux_left_track_167 (
		.in({chany_top_in[141], chany_bottom_in[109], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_60_sram_inv[0:3]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_size12 mux_left_track_169 (
		.in({chany_top_in[140], chany_bottom_in[110], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_61_sram_inv[0:3]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size12 mux_left_track_171 (
		.in({chany_top_in[138], chany_bottom_in[112], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_62_sram_inv[0:3]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_size12 mux_left_track_175 (
		.in({chany_top_in[136], chany_bottom_in[114], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_63_sram_inv[0:3]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_size12 mux_left_track_181 (
		.in({chany_top_in[132], chany_bottom_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_64_sram_inv[0:3]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_size12 mux_left_track_183 (
		.in({chany_top_in[130], chany_bottom_in[120], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_65_sram_inv[0:3]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_size12 mux_left_track_185 (
		.in({chany_top_in[129], chany_bottom_in[121], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_66_sram_inv[0:3]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size12 mux_left_track_187 (
		.in({chany_top_in[128], chany_bottom_in[122], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_67_sram_inv[0:3]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_size12 mux_left_track_189 (
		.in({chany_top_in[126], chany_bottom_in[124], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_68_sram_inv[0:3]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_size12 mux_left_track_191 (
		.in({chany_top_in[125], chany_bottom_in[125], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_69_sram_inv[0:3]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_size12 mux_left_track_199 (
		.in({chany_top_in[120], chany_bottom_in[130], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_70_sram_inv[0:3]),
		.out(chanx_left_out[99]));

	mux_tree_tapbuf_size12 mux_left_track_201 (
		.in({chany_top_in[118], chany_bottom_in[132], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_71_sram_inv[0:3]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size12 mux_left_track_203 (
		.in({chany_top_in[117], chany_bottom_in[133], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_72_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_72_sram_inv[0:3]),
		.out(chanx_left_out[101]));

	mux_tree_tapbuf_size12 mux_left_track_205 (
		.in({chany_top_in[116], chany_bottom_in[134], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_73_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_73_sram_inv[0:3]),
		.out(chanx_left_out[102]));

	mux_tree_tapbuf_size12 mux_left_track_207 (
		.in({chany_top_in[114], chany_bottom_in[136], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_74_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_74_sram_inv[0:3]),
		.out(chanx_left_out[103]));

	mux_tree_tapbuf_size12 mux_left_track_209 (
		.in({chany_top_in[113], chany_bottom_in[137], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_75_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_75_sram_inv[0:3]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size12 mux_left_track_211 (
		.in({chany_top_in[112], chany_bottom_in[138], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_76_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_76_sram_inv[0:3]),
		.out(chanx_left_out[105]));

	mux_tree_tapbuf_size12 mux_left_track_217 (
		.in({chany_top_in[108], chany_bottom_in[142], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_77_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_77_sram_inv[0:3]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size12 mux_left_track_219 (
		.in({chany_top_in[106], chany_bottom_in[144], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_78_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_78_sram_inv[0:3]),
		.out(chanx_left_out[109]));

	mux_tree_tapbuf_size12 mux_left_track_221 (
		.in({chany_top_in[105], chany_bottom_in[145], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_79_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_79_sram_inv[0:3]),
		.out(chanx_left_out[110]));

	mux_tree_tapbuf_size12 mux_left_track_223 (
		.in({chany_top_in[104], chany_bottom_in[146], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_80_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_80_sram_inv[0:3]),
		.out(chanx_left_out[111]));

	mux_tree_tapbuf_size12 mux_left_track_225 (
		.in({chany_top_in[102], chany_bottom_in[148], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_81_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_81_sram_inv[0:3]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size12 mux_left_track_227 (
		.in({chany_top_in[101], chany_bottom_in[149], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_82_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_82_sram_inv[0:3]),
		.out(chanx_left_out[113]));

	mux_tree_tapbuf_size12 mux_left_track_229 (
		.in({chany_top_in[100], chany_bottom_in[150], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_83_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_83_sram_inv[0:3]),
		.out(chanx_left_out[114]));

	mux_tree_tapbuf_size12 mux_left_track_235 (
		.in({chany_top_in[96], chany_bottom_in[154], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_84_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_84_sram_inv[0:3]),
		.out(chanx_left_out[117]));

	mux_tree_tapbuf_size12 mux_left_track_237 (
		.in({chany_top_in[94], chany_bottom_in[156], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_85_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_85_sram_inv[0:3]),
		.out(chanx_left_out[118]));

	mux_tree_tapbuf_size12 mux_left_track_239 (
		.in({chany_top_in[93], chany_bottom_in[157], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_86_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_86_sram_inv[0:3]),
		.out(chanx_left_out[119]));

	mux_tree_tapbuf_size12 mux_left_track_241 (
		.in({chany_top_in[92], chany_bottom_in[158], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_87_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_87_sram_inv[0:3]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size12 mux_left_track_243 (
		.in({chany_top_in[90], chany_bottom_in[160], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_88_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_88_sram_inv[0:3]),
		.out(chanx_left_out[121]));

	mux_tree_tapbuf_size12 mux_left_track_245 (
		.in({chany_top_in[89], chany_bottom_in[161], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_89_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_89_sram_inv[0:3]),
		.out(chanx_left_out[122]));

	mux_tree_tapbuf_size12 mux_left_track_247 (
		.in({chany_top_in[88], chany_bottom_in[162], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_90_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_90_sram_inv[0:3]),
		.out(chanx_left_out[123]));

	mux_tree_tapbuf_size12 mux_left_track_255 (
		.in({chany_top_in[82], chany_bottom_in[168], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_91_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_91_sram_inv[0:3]),
		.out(chanx_left_out[127]));

	mux_tree_tapbuf_size12 mux_left_track_257 (
		.in({chany_top_in[81], chany_bottom_in[169], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_92_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_92_sram_inv[0:3]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size12 mux_left_track_259 (
		.in({chany_top_in[80], chany_bottom_in[170], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_93_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_93_sram_inv[0:3]),
		.out(chanx_left_out[129]));

	mux_tree_tapbuf_size12 mux_left_track_261 (
		.in({chany_top_in[78], chany_bottom_in[172], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_94_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_94_sram_inv[0:3]),
		.out(chanx_left_out[130]));

	mux_tree_tapbuf_size12 mux_left_track_263 (
		.in({chany_top_in[77], chany_bottom_in[173], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_95_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_95_sram_inv[0:3]),
		.out(chanx_left_out[131]));

	mux_tree_tapbuf_size12 mux_left_track_265 (
		.in({chany_top_in[76], chany_bottom_in[174], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_96_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_96_sram_inv[0:3]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size12 mux_left_track_271 (
		.in({chany_top_in[72], chany_bottom_in[178], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_97_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_97_sram_inv[0:3]),
		.out(chanx_left_out[135]));

	mux_tree_tapbuf_size12 mux_left_track_275 (
		.in({chany_top_in[69], chany_bottom_in[181], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_98_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_98_sram_inv[0:3]),
		.out(chanx_left_out[137]));

	mux_tree_tapbuf_size12 mux_left_track_277 (
		.in({chany_top_in[68], chany_bottom_in[182], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_99_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_99_sram_inv[0:3]),
		.out(chanx_left_out[138]));

	mux_tree_tapbuf_size12 mux_left_track_279 (
		.in({chany_top_in[66], chany_bottom_in[184], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size12_100_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_100_sram_inv[0:3]),
		.out(chanx_left_out[139]));

	mux_tree_tapbuf_size12 mux_left_track_281 (
		.in({chany_top_in[65], chany_bottom_in[185], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_101_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_101_sram_inv[0:3]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size12 mux_left_track_283 (
		.in({chany_top_in[64], chany_bottom_in[186], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_102_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_102_sram_inv[0:3]),
		.out(chanx_left_out[141]));

	mux_tree_tapbuf_size12 mux_left_track_289 (
		.in({chany_top_in[60], chany_top_in[183], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_103_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_103_sram_inv[0:3]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size12 mux_left_track_291 (
		.in({chany_top_in[58], chany_top_in[179], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_104_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_104_sram_inv[0:3]),
		.out(chanx_left_out[145]));

	mux_tree_tapbuf_size12 mux_left_track_295 (
		.in({chany_top_in[56], chany_top_in[171], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_105_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_105_sram_inv[0:3]),
		.out(chanx_left_out[147]));

	mux_tree_tapbuf_size12 mux_left_track_297 (
		.in({chany_top_in[54], chany_top_in[167], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_106_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_106_sram_inv[0:3]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size12 mux_left_track_299 (
		.in({chany_top_in[53], chany_top_in[163], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_107_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_107_sram_inv[0:3]),
		.out(chanx_left_out[149]));

	mux_tree_tapbuf_size12 mux_left_track_301 (
		.in({chany_top_in[52], chany_top_in[159], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_108_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_108_sram_inv[0:3]),
		.out(chanx_left_out[150]));

	mux_tree_tapbuf_size12 mux_left_track_307 (
		.in({chany_top_in[48], chany_top_in[147], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_109_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_109_sram_inv[0:3]),
		.out(chanx_left_out[153]));

	mux_tree_tapbuf_size12 mux_left_track_309 (
		.in({chany_top_in[46], chany_top_in[143], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_110_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_110_sram_inv[0:3]),
		.out(chanx_left_out[154]));

	mux_tree_tapbuf_size12 mux_left_track_311 (
		.in({chany_top_in[45], chany_top_in[139], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_111_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_111_sram_inv[0:3]),
		.out(chanx_left_out[155]));

	mux_tree_tapbuf_size12 mux_left_track_315 (
		.in({chany_top_in[42], chany_top_in[131], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size12_112_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_112_sram_inv[0:3]),
		.out(chanx_left_out[157]));

	mux_tree_tapbuf_size12 mux_left_track_317 (
		.in({chany_top_in[41], chany_top_in[127], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_113_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_113_sram_inv[0:3]),
		.out(chanx_left_out[158]));

	mux_tree_tapbuf_size12 mux_left_track_319 (
		.in({chany_top_in[40], chany_top_in[123], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_114_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_114_sram_inv[0:3]),
		.out(chanx_left_out[159]));

	mux_tree_tapbuf_size12 mux_left_track_325 (
		.in({chany_top_in[36], chany_top_in[111], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_115_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_115_sram_inv[0:3]),
		.out(chanx_left_out[162]));

	mux_tree_tapbuf_size12 mux_left_track_327 (
		.in({chany_top_in[34], chany_top_in[107], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_116_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_116_sram_inv[0:3]),
		.out(chanx_left_out[163]));

	mux_tree_tapbuf_size12 mux_left_track_329 (
		.in({chany_top_in[33], chany_top_in[103], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_117_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_117_sram_inv[0:3]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size12 mux_left_track_331 (
		.in({chany_top_in[32], chany_top_in[99], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_118_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_118_sram_inv[0:3]),
		.out(chanx_left_out[165]));

	mux_tree_tapbuf_size12 mux_left_track_335 (
		.in({chany_top_in[29], chany_top_in[91], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_119_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_119_sram_inv[0:3]),
		.out(chanx_left_out[167]));

	mux_tree_tapbuf_size12 mux_left_track_337 (
		.in({chany_top_in[28], chany_top_in[87], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_120_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_120_sram_inv[0:3]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size12 mux_left_track_343 (
		.in({chany_top_in[24], chany_top_in[75], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_121_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_121_sram_inv[0:3]),
		.out(chanx_left_out[171]));

	mux_tree_tapbuf_size12 mux_left_track_345 (
		.in({chany_top_in[22], chany_top_in[71], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_122_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_122_sram_inv[0:3]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size12 mux_left_track_347 (
		.in({chany_top_in[21], chany_top_in[67], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_123_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_123_sram_inv[0:3]),
		.out(chanx_left_out[173]));

	mux_tree_tapbuf_size12 mux_left_track_349 (
		.in({chany_top_in[20], chany_top_in[63], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_124_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_124_sram_inv[0:3]),
		.out(chanx_left_out[174]));

	mux_tree_tapbuf_size12 mux_left_track_351 (
		.in({chany_top_in[18], chany_top_in[59], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size12_125_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_125_sram_inv[0:3]),
		.out(chanx_left_out[175]));

	mux_tree_tapbuf_size12 mux_left_track_355 (
		.in({chany_top_in[16], chany_top_in[51], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size12_126_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_126_sram_inv[0:3]),
		.out(chanx_left_out[177]));

	mux_tree_tapbuf_size12 mux_left_track_361 (
		.in({chany_top_in[12], chany_top_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size12_127_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_127_sram_inv[0:3]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size12 mux_left_track_363 (
		.in({chany_top_in[10], chany_top_in[35], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size12_128_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_128_sram_inv[0:3]),
		.out(chanx_left_out[181]));

	mux_tree_tapbuf_size12 mux_left_track_365 (
		.in({chany_top_in[9], chany_top_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size12_129_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_129_sram_inv[0:3]),
		.out(chanx_left_out[182]));

	mux_tree_tapbuf_size12 mux_left_track_367 (
		.in({chany_top_in[8], chany_top_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_130_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_130_sram_inv[0:3]),
		.out(chanx_left_out[183]));

	mux_tree_tapbuf_size12 mux_left_track_369 (
		.in({chany_top_in[6], chany_top_in[23], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_131_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_131_sram_inv[0:3]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size12 mux_left_track_371 (
		.in({chany_top_in[5], chany_top_in[19], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size12_132_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_132_sram_inv[0:3]),
		.out(chanx_left_out[185]));

	mux_tree_tapbuf_size12_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size16_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_36_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_37_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_38_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_39_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_40_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_41_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_42_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_43_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_44_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_45_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_46_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_47_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_48_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_49_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_50_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_51_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_52_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_53_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_54_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_55_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_56_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_57_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_58_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_59_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_60_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_61_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_62_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_63_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_64_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_65_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_66_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_67_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_68_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_69_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_70_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_71_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_72_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_72_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_73_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_73_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_74_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_74_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_75_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_75_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_76_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_76_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_77_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_77_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_219 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_78_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_78_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_221 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_79_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_79_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_223 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_80_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_80_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_81_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_81_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_227 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_82_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_82_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_229 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_83_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_83_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_235 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_84_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_84_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_237 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_85_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_85_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_239 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_86_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_86_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_87_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_87_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_243 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_88_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_88_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_245 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_89_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_89_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_247 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_90_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_90_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_255 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_91_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_91_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_92_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_92_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_259 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_93_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_93_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_261 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_94_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_94_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_263 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_95_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_95_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_96_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_96_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_271 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_97_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_97_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_275 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_98_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_98_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_277 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_99_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_99_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_279 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_100_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_100_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_101_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_101_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_283 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_102_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_102_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_103_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_103_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_291 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_104_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_104_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_295 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_105_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_105_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_106_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_106_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_299 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_107_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_107_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_301 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_108_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_108_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_307 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_109_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_109_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_309 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_110_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_110_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_311 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_111_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_111_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_315 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_112_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_112_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_317 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_113_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_113_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_319 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_114_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_114_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_325 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_115_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_115_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_327 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_116_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_116_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_117_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_117_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_331 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_118_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_118_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_335 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_119_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_119_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_120_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_120_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_343 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_121_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_121_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_122_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_122_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_347 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_123_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_123_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_349 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_124_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_124_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_351 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_125_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_125_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_355 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_126_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_126_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_127_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_127_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_363 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_128_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_128_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_365 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_129_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_129_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_367 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_130_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_130_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_131_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_131_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_left_track_371 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_132_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_132_sram_inv[0:3]));

	mux_tree_tapbuf_size10 mux_left_track_15 (
		.in({chany_bottom_in[8], chany_bottom_in[27], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size10 mux_left_track_35 (
		.in({chany_bottom_in[21], chany_bottom_in[67], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_}),
		.sram(mux_tree_tapbuf_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_1_sram_inv[0:3]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size10 mux_left_track_213 (
		.in({chany_top_in[110], chany_bottom_in[140], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_}),
		.sram(mux_tree_tapbuf_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_2_sram_inv[0:3]),
		.out(chanx_left_out[106]));

	mux_tree_tapbuf_size10 mux_left_track_233 (
		.in({chany_top_in[97], chany_bottom_in[153], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_}),
		.sram(mux_tree_tapbuf_size10_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_3_sram_inv[0:3]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size10_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_213 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11 mux_left_track_17 (
		.in({chany_bottom_in[9], chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size11 mux_left_track_33 (
		.in({chany_bottom_in[20], chany_bottom_in[63], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size11 mux_left_track_51 (
		.in({chany_bottom_in[32], chany_bottom_in[99], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size11 mux_left_track_53 (
		.in({chany_bottom_in[33], chany_bottom_in[103], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size11 mux_left_track_55 (
		.in({chany_bottom_in[34], chany_bottom_in[107], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size11 mux_left_track_69 (
		.in({chany_bottom_in[44], chany_bottom_in[135], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size11 mux_left_track_71 (
		.in({chany_bottom_in[45], chany_bottom_in[139], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size11 mux_left_track_75 (
		.in({chany_bottom_in[48], chany_bottom_in[147], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size11 mux_left_track_87 (
		.in({chany_bottom_in[56], chany_bottom_in[171], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size11 mux_left_track_89 (
		.in({chany_bottom_in[57], chany_bottom_in[175], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size11 mux_left_track_95 (
		.in({chany_bottom_in[61], chany_bottom_in[187], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size11 mux_left_track_105 (
		.in({chany_top_in[182], chany_bottom_in[68], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_11_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size11 mux_left_track_107 (
		.in({chany_top_in[181], chany_bottom_in[69], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_12_sram_inv[0:3]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size11 mux_left_track_115 (
		.in({chany_top_in[176], chany_bottom_in[74], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_}),
		.sram(mux_tree_tapbuf_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_13_sram_inv[0:3]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size11 mux_left_track_123 (
		.in({chany_top_in[170], chany_bottom_in[80], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_14_sram_inv[0:3]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size11 mux_left_track_125 (
		.in({chany_top_in[169], chany_bottom_in[81], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size11_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_15_sram_inv[0:3]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size11 mux_left_track_135 (
		.in({chany_top_in[162], chany_bottom_in[88], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size11_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_16_sram_inv[0:3]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size11 mux_left_track_141 (
		.in({chany_top_in[158], chany_bottom_in[92], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_17_sram_inv[0:3]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size11 mux_left_track_143 (
		.in({chany_top_in[157], chany_bottom_in[93], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_18_sram_inv[0:3]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size11 mux_left_track_159 (
		.in({chany_top_in[146], chany_bottom_in[104], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_19_sram_inv[0:3]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_size11 mux_left_track_161 (
		.in({chany_top_in[145], chany_bottom_in[105], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_20_sram_inv[0:3]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size11 mux_left_track_173 (
		.in({chany_top_in[137], chany_bottom_in[113], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size11_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_21_sram_inv[0:3]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_size11 mux_left_track_177 (
		.in({chany_top_in[134], chany_bottom_in[116], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_22_sram_inv[0:3]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size11 mux_left_track_179 (
		.in({chany_top_in[133], chany_bottom_in[117], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_23_sram_inv[0:3]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_size11 mux_left_track_193 (
		.in({chany_top_in[124], chany_bottom_in[126], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size11_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_24_sram_inv[0:3]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size11 mux_left_track_195 (
		.in({chany_top_in[122], chany_bottom_in[128], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size11_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_25_sram_inv[0:3]),
		.out(chanx_left_out[97]));

	mux_tree_tapbuf_size11 mux_left_track_197 (
		.in({chany_top_in[121], chany_bottom_in[129], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_26_sram_inv[0:3]),
		.out(chanx_left_out[98]));

	mux_tree_tapbuf_size11 mux_left_track_215 (
		.in({chany_top_in[109], chany_bottom_in[141], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size11_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_27_sram_inv[0:3]),
		.out(chanx_left_out[107]));

	mux_tree_tapbuf_size11 mux_left_track_231 (
		.in({chany_top_in[98], chany_bottom_in[152], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size11_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_28_sram_inv[0:3]),
		.out(chanx_left_out[115]));

	mux_tree_tapbuf_size11 mux_left_track_249 (
		.in({chany_top_in[86], chany_bottom_in[164], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size11_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_29_sram_inv[0:3]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size11 mux_left_track_251 (
		.in({chany_top_in[85], chany_bottom_in[165], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size11_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_30_sram_inv[0:3]),
		.out(chanx_left_out[125]));

	mux_tree_tapbuf_size11 mux_left_track_253 (
		.in({chany_top_in[84], chany_bottom_in[166], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_}),
		.sram(mux_tree_tapbuf_size11_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_31_sram_inv[0:3]),
		.out(chanx_left_out[126]));

	mux_tree_tapbuf_size11 mux_left_track_267 (
		.in({chany_top_in[74], chany_bottom_in[176], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size11_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_32_sram_inv[0:3]),
		.out(chanx_left_out[133]));

	mux_tree_tapbuf_size11 mux_left_track_269 (
		.in({chany_top_in[73], chany_bottom_in[177], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size11_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_33_sram_inv[0:3]),
		.out(chanx_left_out[134]));

	mux_tree_tapbuf_size11 mux_left_track_273 (
		.in({chany_top_in[70], chany_bottom_in[180], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_}),
		.sram(mux_tree_tapbuf_size11_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_34_sram_inv[0:3]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size11 mux_left_track_285 (
		.in({chany_top_in[62], chany_top_in[188], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size11_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_35_sram_inv[0:3]),
		.out(chanx_left_out[142]));

	mux_tree_tapbuf_size11 mux_left_track_287 (
		.in({chany_top_in[61], chany_top_in[187], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size11_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_36_sram_inv[0:3]),
		.out(chanx_left_out[143]));

	mux_tree_tapbuf_size11 mux_left_track_293 (
		.in({chany_top_in[57], chany_top_in[175], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_}),
		.sram(mux_tree_tapbuf_size11_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_37_sram_inv[0:3]),
		.out(chanx_left_out[146]));

	mux_tree_tapbuf_size11 mux_left_track_303 (
		.in({chany_top_in[50], chany_top_in[155], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size11_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_38_sram_inv[0:3]),
		.out(chanx_left_out[151]));

	mux_tree_tapbuf_size11 mux_left_track_305 (
		.in({chany_top_in[49], chany_top_in[151], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size11_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_39_sram_inv[0:3]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size11 mux_left_track_313 (
		.in({chany_top_in[44], chany_top_in[135], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_}),
		.sram(mux_tree_tapbuf_size11_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_40_sram_inv[0:3]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size11 mux_left_track_321 (
		.in({chany_top_in[38], chany_top_in[119], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_41_sram_inv[0:3]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size11 mux_left_track_323 (
		.in({chany_top_in[37], chany_top_in[115], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size11_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_42_sram_inv[0:3]),
		.out(chanx_left_out[161]));

	mux_tree_tapbuf_size11 mux_left_track_333 (
		.in({chany_top_in[30], chany_top_in[95], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size11_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_43_sram_inv[0:3]),
		.out(chanx_left_out[166]));

	mux_tree_tapbuf_size11 mux_left_track_339 (
		.in({chany_top_in[26], chany_top_in[83], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_44_sram_inv[0:3]),
		.out(chanx_left_out[169]));

	mux_tree_tapbuf_size11 mux_left_track_341 (
		.in({chany_top_in[25], chany_top_in[79], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_45_sram_inv[0:3]),
		.out(chanx_left_out[170]));

	mux_tree_tapbuf_size11 mux_left_track_353 (
		.in({chany_top_in[17], chany_top_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size11_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_46_sram_inv[0:3]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size11 mux_left_track_357 (
		.in({chany_top_in[14], chany_top_in[47], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_47_sram_inv[0:3]),
		.out(chanx_left_out[178]));

	mux_tree_tapbuf_size11 mux_left_track_359 (
		.in({chany_top_in[13], chany_top_in[43], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_48_sram_inv[0:3]),
		.out(chanx_left_out[179]));

	mux_tree_tapbuf_size11 mux_left_track_373 (
		.in({chany_top_in[4], chany_top_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size11_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_49_sram_inv[0:3]),
		.out(chanx_left_out[186]));

	mux_tree_tapbuf_size11 mux_left_track_375 (
		.in({chany_top_in[2], chany_top_in[11], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_}),
		.sram(mux_tree_tapbuf_size11_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_50_sram_inv[0:3]),
		.out(chanx_left_out[187]));

	mux_tree_tapbuf_size11 mux_left_track_377 (
		.in({chany_top_in[1], chany_top_in[7], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size11_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_51_sram_inv[0:3]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size11_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_14_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_15_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_16_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_17_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_18_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_19_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_20_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_21_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_22_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_23_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_24_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_25_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_26_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_215 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_27_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_231 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_28_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_29_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_251 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_30_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_253 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_31_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_267 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_32_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_269 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_33_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_34_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_285 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_35_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_287 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_36_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_293 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_37_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_303 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_38_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_39_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_40_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_41_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_323 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_42_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_333 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_43_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_339 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_44_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_341 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_45_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_46_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_357 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_47_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_359 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_48_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_373 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_49_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_375 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_50_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_50_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_51_sram_inv[0:3]));

endmodule
// ----- END Verilog module for sb_4__2_ -----

//----- Default net type -----
`default_nettype wire



