//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Formal Top-level netlist of Design: router_mesh
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul  7 02:20:28 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module router_mesh_top_formal_verification_random_tb;
// ----- Default clock port is added here since benchmark does not contain one -------
	reg [0:0] clk;

// ----- Shared inputs -------
	reg [0:0] reset;
	reg [0:0] injection_channels_629_;
	reg [0:0] injection_channels_628_;
	reg [0:0] injection_channels_627_;
	reg [0:0] injection_channels_626_;
	reg [0:0] injection_channels_625_;
	reg [0:0] injection_channels_624_;
	reg [0:0] injection_channels_623_;
	reg [0:0] injection_channels_622_;
	reg [0:0] injection_channels_621_;
	reg [0:0] injection_channels_620_;
	reg [0:0] injection_channels_619_;
	reg [0:0] injection_channels_618_;
	reg [0:0] injection_channels_617_;
	reg [0:0] injection_channels_616_;
	reg [0:0] injection_channels_615_;
	reg [0:0] injection_channels_614_;
	reg [0:0] injection_channels_613_;
	reg [0:0] injection_channels_612_;
	reg [0:0] injection_channels_611_;
	reg [0:0] injection_channels_610_;
	reg [0:0] injection_channels_609_;
	reg [0:0] injection_channels_608_;
	reg [0:0] injection_channels_607_;
	reg [0:0] injection_channels_606_;
	reg [0:0] injection_channels_605_;
	reg [0:0] injection_channels_604_;
	reg [0:0] injection_channels_603_;
	reg [0:0] injection_channels_602_;
	reg [0:0] injection_channels_601_;
	reg [0:0] injection_channels_600_;
	reg [0:0] injection_channels_599_;
	reg [0:0] injection_channels_598_;
	reg [0:0] injection_channels_597_;
	reg [0:0] injection_channels_596_;
	reg [0:0] injection_channels_595_;
	reg [0:0] injection_channels_594_;
	reg [0:0] injection_channels_593_;
	reg [0:0] injection_channels_592_;
	reg [0:0] injection_channels_591_;
	reg [0:0] injection_channels_590_;
	reg [0:0] injection_channels_589_;
	reg [0:0] injection_channels_588_;
	reg [0:0] injection_channels_587_;
	reg [0:0] injection_channels_586_;
	reg [0:0] injection_channels_585_;
	reg [0:0] injection_channels_584_;
	reg [0:0] injection_channels_583_;
	reg [0:0] injection_channels_582_;
	reg [0:0] injection_channels_581_;
	reg [0:0] injection_channels_580_;
	reg [0:0] injection_channels_579_;
	reg [0:0] injection_channels_578_;
	reg [0:0] injection_channels_577_;
	reg [0:0] injection_channels_576_;
	reg [0:0] injection_channels_575_;
	reg [0:0] injection_channels_574_;
	reg [0:0] injection_channels_573_;
	reg [0:0] injection_channels_572_;
	reg [0:0] injection_channels_571_;
	reg [0:0] injection_channels_570_;
	reg [0:0] injection_channels_569_;
	reg [0:0] injection_channels_568_;
	reg [0:0] injection_channels_567_;
	reg [0:0] injection_channels_566_;
	reg [0:0] injection_channels_565_;
	reg [0:0] injection_channels_564_;
	reg [0:0] injection_channels_563_;
	reg [0:0] injection_channels_562_;
	reg [0:0] injection_channels_561_;
	reg [0:0] injection_channels_560_;
	reg [0:0] injection_channels_559_;
	reg [0:0] injection_channels_558_;
	reg [0:0] injection_channels_557_;
	reg [0:0] injection_channels_556_;
	reg [0:0] injection_channels_555_;
	reg [0:0] injection_channels_554_;
	reg [0:0] injection_channels_553_;
	reg [0:0] injection_channels_552_;
	reg [0:0] injection_channels_551_;
	reg [0:0] injection_channels_550_;
	reg [0:0] injection_channels_549_;
	reg [0:0] injection_channels_548_;
	reg [0:0] injection_channels_547_;
	reg [0:0] injection_channels_546_;
	reg [0:0] injection_channels_545_;
	reg [0:0] injection_channels_544_;
	reg [0:0] injection_channels_543_;
	reg [0:0] injection_channels_542_;
	reg [0:0] injection_channels_541_;
	reg [0:0] injection_channels_540_;
	reg [0:0] injection_channels_539_;
	reg [0:0] injection_channels_538_;
	reg [0:0] injection_channels_537_;
	reg [0:0] injection_channels_536_;
	reg [0:0] injection_channels_535_;
	reg [0:0] injection_channels_534_;
	reg [0:0] injection_channels_533_;
	reg [0:0] injection_channels_532_;
	reg [0:0] injection_channels_531_;
	reg [0:0] injection_channels_530_;
	reg [0:0] injection_channels_529_;
	reg [0:0] injection_channels_528_;
	reg [0:0] injection_channels_527_;
	reg [0:0] injection_channels_526_;
	reg [0:0] injection_channels_525_;
	reg [0:0] injection_channels_524_;
	reg [0:0] injection_channels_523_;
	reg [0:0] injection_channels_522_;
	reg [0:0] injection_channels_521_;
	reg [0:0] injection_channels_520_;
	reg [0:0] injection_channels_519_;
	reg [0:0] injection_channels_518_;
	reg [0:0] injection_channels_517_;
	reg [0:0] injection_channels_516_;
	reg [0:0] injection_channels_515_;
	reg [0:0] injection_channels_514_;
	reg [0:0] injection_channels_513_;
	reg [0:0] injection_channels_512_;
	reg [0:0] injection_channels_511_;
	reg [0:0] injection_channels_510_;
	reg [0:0] injection_channels_509_;
	reg [0:0] injection_channels_508_;
	reg [0:0] injection_channels_507_;
	reg [0:0] injection_channels_506_;
	reg [0:0] injection_channels_505_;
	reg [0:0] injection_channels_504_;
	reg [0:0] injection_channels_503_;
	reg [0:0] injection_channels_502_;
	reg [0:0] injection_channels_501_;
	reg [0:0] injection_channels_500_;
	reg [0:0] injection_channels_499_;
	reg [0:0] injection_channels_498_;
	reg [0:0] injection_channels_497_;
	reg [0:0] injection_channels_496_;
	reg [0:0] injection_channels_495_;
	reg [0:0] injection_channels_494_;
	reg [0:0] injection_channels_493_;
	reg [0:0] injection_channels_492_;
	reg [0:0] injection_channels_491_;
	reg [0:0] injection_channels_490_;
	reg [0:0] injection_channels_489_;
	reg [0:0] injection_channels_488_;
	reg [0:0] injection_channels_487_;
	reg [0:0] injection_channels_486_;
	reg [0:0] injection_channels_485_;
	reg [0:0] injection_channels_484_;
	reg [0:0] injection_channels_483_;
	reg [0:0] injection_channels_482_;
	reg [0:0] injection_channels_481_;
	reg [0:0] injection_channels_480_;
	reg [0:0] injection_channels_479_;
	reg [0:0] injection_channels_478_;
	reg [0:0] injection_channels_477_;
	reg [0:0] injection_channels_476_;
	reg [0:0] injection_channels_475_;
	reg [0:0] injection_channels_474_;
	reg [0:0] injection_channels_473_;
	reg [0:0] injection_channels_472_;
	reg [0:0] injection_channels_471_;
	reg [0:0] injection_channels_470_;
	reg [0:0] injection_channels_469_;
	reg [0:0] injection_channels_468_;
	reg [0:0] injection_channels_467_;
	reg [0:0] injection_channels_466_;
	reg [0:0] injection_channels_465_;
	reg [0:0] injection_channels_464_;
	reg [0:0] injection_channels_463_;
	reg [0:0] injection_channels_462_;
	reg [0:0] injection_channels_461_;
	reg [0:0] injection_channels_460_;
	reg [0:0] injection_channels_459_;
	reg [0:0] injection_channels_458_;
	reg [0:0] injection_channels_457_;
	reg [0:0] injection_channels_456_;
	reg [0:0] injection_channels_455_;
	reg [0:0] injection_channels_454_;
	reg [0:0] injection_channels_453_;
	reg [0:0] injection_channels_452_;
	reg [0:0] injection_channels_451_;
	reg [0:0] injection_channels_450_;
	reg [0:0] injection_channels_449_;
	reg [0:0] injection_channels_448_;
	reg [0:0] injection_channels_447_;
	reg [0:0] injection_channels_446_;
	reg [0:0] injection_channels_445_;
	reg [0:0] injection_channels_444_;
	reg [0:0] injection_channels_443_;
	reg [0:0] injection_channels_442_;
	reg [0:0] injection_channels_441_;
	reg [0:0] injection_channels_440_;
	reg [0:0] injection_channels_439_;
	reg [0:0] injection_channels_438_;
	reg [0:0] injection_channels_437_;
	reg [0:0] injection_channels_436_;
	reg [0:0] injection_channels_435_;
	reg [0:0] injection_channels_434_;
	reg [0:0] injection_channels_433_;
	reg [0:0] injection_channels_432_;
	reg [0:0] injection_channels_431_;
	reg [0:0] injection_channels_430_;
	reg [0:0] injection_channels_429_;
	reg [0:0] injection_channels_428_;
	reg [0:0] injection_channels_427_;
	reg [0:0] injection_channels_426_;
	reg [0:0] injection_channels_425_;
	reg [0:0] injection_channels_424_;
	reg [0:0] injection_channels_423_;
	reg [0:0] injection_channels_422_;
	reg [0:0] injection_channels_421_;
	reg [0:0] injection_channels_420_;
	reg [0:0] injection_channels_419_;
	reg [0:0] injection_channels_418_;
	reg [0:0] injection_channels_417_;
	reg [0:0] injection_channels_416_;
	reg [0:0] injection_channels_415_;
	reg [0:0] injection_channels_414_;
	reg [0:0] injection_channels_413_;
	reg [0:0] injection_channels_412_;
	reg [0:0] injection_channels_411_;
	reg [0:0] injection_channels_410_;
	reg [0:0] injection_channels_409_;
	reg [0:0] injection_channels_408_;
	reg [0:0] injection_channels_407_;
	reg [0:0] injection_channels_406_;
	reg [0:0] injection_channels_405_;
	reg [0:0] injection_channels_404_;
	reg [0:0] injection_channels_403_;
	reg [0:0] injection_channels_402_;
	reg [0:0] injection_channels_401_;
	reg [0:0] injection_channels_400_;
	reg [0:0] injection_channels_399_;
	reg [0:0] injection_channels_398_;
	reg [0:0] injection_channels_397_;
	reg [0:0] injection_channels_396_;
	reg [0:0] injection_channels_395_;
	reg [0:0] injection_channels_394_;
	reg [0:0] injection_channels_393_;
	reg [0:0] injection_channels_392_;
	reg [0:0] injection_channels_391_;
	reg [0:0] injection_channels_390_;
	reg [0:0] injection_channels_389_;
	reg [0:0] injection_channels_388_;
	reg [0:0] injection_channels_387_;
	reg [0:0] injection_channels_386_;
	reg [0:0] injection_channels_385_;
	reg [0:0] injection_channels_384_;
	reg [0:0] injection_channels_383_;
	reg [0:0] injection_channels_382_;
	reg [0:0] injection_channels_381_;
	reg [0:0] injection_channels_380_;
	reg [0:0] injection_channels_379_;
	reg [0:0] injection_channels_378_;
	reg [0:0] injection_channels_377_;
	reg [0:0] injection_channels_376_;
	reg [0:0] injection_channels_375_;
	reg [0:0] injection_channels_374_;
	reg [0:0] injection_channels_373_;
	reg [0:0] injection_channels_372_;
	reg [0:0] injection_channels_371_;
	reg [0:0] injection_channels_370_;
	reg [0:0] injection_channels_369_;
	reg [0:0] injection_channels_368_;
	reg [0:0] injection_channels_367_;
	reg [0:0] injection_channels_366_;
	reg [0:0] injection_channels_365_;
	reg [0:0] injection_channels_364_;
	reg [0:0] injection_channels_363_;
	reg [0:0] injection_channels_362_;
	reg [0:0] injection_channels_361_;
	reg [0:0] injection_channels_360_;
	reg [0:0] injection_channels_359_;
	reg [0:0] injection_channels_358_;
	reg [0:0] injection_channels_357_;
	reg [0:0] injection_channels_356_;
	reg [0:0] injection_channels_355_;
	reg [0:0] injection_channels_354_;
	reg [0:0] injection_channels_353_;
	reg [0:0] injection_channels_352_;
	reg [0:0] injection_channels_351_;
	reg [0:0] injection_channels_350_;
	reg [0:0] injection_channels_349_;
	reg [0:0] injection_channels_348_;
	reg [0:0] injection_channels_347_;
	reg [0:0] injection_channels_346_;
	reg [0:0] injection_channels_345_;
	reg [0:0] injection_channels_344_;
	reg [0:0] injection_channels_343_;
	reg [0:0] injection_channels_342_;
	reg [0:0] injection_channels_341_;
	reg [0:0] injection_channels_340_;
	reg [0:0] injection_channels_339_;
	reg [0:0] injection_channels_338_;
	reg [0:0] injection_channels_337_;
	reg [0:0] injection_channels_336_;
	reg [0:0] injection_channels_335_;
	reg [0:0] injection_channels_334_;
	reg [0:0] injection_channels_333_;
	reg [0:0] injection_channels_332_;
	reg [0:0] injection_channels_331_;
	reg [0:0] injection_channels_330_;
	reg [0:0] injection_channels_329_;
	reg [0:0] injection_channels_328_;
	reg [0:0] injection_channels_327_;
	reg [0:0] injection_channels_326_;
	reg [0:0] injection_channels_325_;
	reg [0:0] injection_channels_324_;
	reg [0:0] injection_channels_323_;
	reg [0:0] injection_channels_322_;
	reg [0:0] injection_channels_321_;
	reg [0:0] injection_channels_320_;
	reg [0:0] injection_channels_319_;
	reg [0:0] injection_channels_318_;
	reg [0:0] injection_channels_317_;
	reg [0:0] injection_channels_316_;
	reg [0:0] injection_channels_315_;
	reg [0:0] injection_channels_314_;
	reg [0:0] injection_channels_313_;
	reg [0:0] injection_channels_312_;
	reg [0:0] injection_channels_311_;
	reg [0:0] injection_channels_310_;
	reg [0:0] injection_channels_309_;
	reg [0:0] injection_channels_308_;
	reg [0:0] injection_channels_307_;
	reg [0:0] injection_channels_306_;
	reg [0:0] injection_channels_305_;
	reg [0:0] injection_channels_304_;
	reg [0:0] injection_channels_303_;
	reg [0:0] injection_channels_302_;
	reg [0:0] injection_channels_301_;
	reg [0:0] injection_channels_300_;
	reg [0:0] injection_channels_299_;
	reg [0:0] injection_channels_298_;
	reg [0:0] injection_channels_297_;
	reg [0:0] injection_channels_296_;
	reg [0:0] injection_channels_295_;
	reg [0:0] injection_channels_294_;
	reg [0:0] injection_channels_293_;
	reg [0:0] injection_channels_292_;
	reg [0:0] injection_channels_291_;
	reg [0:0] injection_channels_290_;
	reg [0:0] injection_channels_289_;
	reg [0:0] injection_channels_288_;
	reg [0:0] injection_channels_287_;
	reg [0:0] injection_channels_286_;
	reg [0:0] injection_channels_285_;
	reg [0:0] injection_channels_284_;
	reg [0:0] injection_channels_283_;
	reg [0:0] injection_channels_282_;
	reg [0:0] injection_channels_281_;
	reg [0:0] injection_channels_280_;
	reg [0:0] injection_channels_279_;
	reg [0:0] injection_channels_278_;
	reg [0:0] injection_channels_277_;
	reg [0:0] injection_channels_276_;
	reg [0:0] injection_channels_275_;
	reg [0:0] injection_channels_274_;
	reg [0:0] injection_channels_273_;
	reg [0:0] injection_channels_272_;
	reg [0:0] injection_channels_271_;
	reg [0:0] injection_channels_270_;
	reg [0:0] injection_channels_269_;
	reg [0:0] injection_channels_268_;
	reg [0:0] injection_channels_267_;
	reg [0:0] injection_channels_266_;
	reg [0:0] injection_channels_265_;
	reg [0:0] injection_channels_264_;
	reg [0:0] injection_channels_263_;
	reg [0:0] injection_channels_262_;
	reg [0:0] injection_channels_261_;
	reg [0:0] injection_channels_260_;
	reg [0:0] injection_channels_259_;
	reg [0:0] injection_channels_258_;
	reg [0:0] injection_channels_257_;
	reg [0:0] injection_channels_256_;
	reg [0:0] injection_channels_255_;
	reg [0:0] injection_channels_254_;
	reg [0:0] injection_channels_253_;
	reg [0:0] injection_channels_252_;
	reg [0:0] injection_channels_251_;
	reg [0:0] injection_channels_250_;
	reg [0:0] injection_channels_249_;
	reg [0:0] injection_channels_248_;
	reg [0:0] injection_channels_247_;
	reg [0:0] injection_channels_246_;
	reg [0:0] injection_channels_245_;
	reg [0:0] injection_channels_244_;
	reg [0:0] injection_channels_243_;
	reg [0:0] injection_channels_242_;
	reg [0:0] injection_channels_241_;
	reg [0:0] injection_channels_240_;
	reg [0:0] injection_channels_239_;
	reg [0:0] injection_channels_238_;
	reg [0:0] injection_channels_237_;
	reg [0:0] injection_channels_236_;
	reg [0:0] injection_channels_235_;
	reg [0:0] injection_channels_234_;
	reg [0:0] injection_channels_233_;
	reg [0:0] injection_channels_232_;
	reg [0:0] injection_channels_231_;
	reg [0:0] injection_channels_230_;
	reg [0:0] injection_channels_229_;
	reg [0:0] injection_channels_228_;
	reg [0:0] injection_channels_227_;
	reg [0:0] injection_channels_226_;
	reg [0:0] injection_channels_225_;
	reg [0:0] injection_channels_224_;
	reg [0:0] injection_channels_223_;
	reg [0:0] injection_channels_222_;
	reg [0:0] injection_channels_221_;
	reg [0:0] injection_channels_220_;
	reg [0:0] injection_channels_219_;
	reg [0:0] injection_channels_218_;
	reg [0:0] injection_channels_217_;
	reg [0:0] injection_channels_216_;
	reg [0:0] injection_channels_215_;
	reg [0:0] injection_channels_214_;
	reg [0:0] injection_channels_213_;
	reg [0:0] injection_channels_212_;
	reg [0:0] injection_channels_211_;
	reg [0:0] injection_channels_210_;
	reg [0:0] injection_channels_209_;
	reg [0:0] injection_channels_208_;
	reg [0:0] injection_channels_207_;
	reg [0:0] injection_channels_206_;
	reg [0:0] injection_channels_205_;
	reg [0:0] injection_channels_204_;
	reg [0:0] injection_channels_203_;
	reg [0:0] injection_channels_202_;
	reg [0:0] injection_channels_201_;
	reg [0:0] injection_channels_200_;
	reg [0:0] injection_channels_199_;
	reg [0:0] injection_channels_198_;
	reg [0:0] injection_channels_197_;
	reg [0:0] injection_channels_196_;
	reg [0:0] injection_channels_195_;
	reg [0:0] injection_channels_194_;
	reg [0:0] injection_channels_193_;
	reg [0:0] injection_channels_192_;
	reg [0:0] injection_channels_191_;
	reg [0:0] injection_channels_190_;
	reg [0:0] injection_channels_189_;
	reg [0:0] injection_channels_188_;
	reg [0:0] injection_channels_187_;
	reg [0:0] injection_channels_186_;
	reg [0:0] injection_channels_185_;
	reg [0:0] injection_channels_184_;
	reg [0:0] injection_channels_183_;
	reg [0:0] injection_channels_182_;
	reg [0:0] injection_channels_181_;
	reg [0:0] injection_channels_180_;
	reg [0:0] injection_channels_179_;
	reg [0:0] injection_channels_178_;
	reg [0:0] injection_channels_177_;
	reg [0:0] injection_channels_176_;
	reg [0:0] injection_channels_175_;
	reg [0:0] injection_channels_174_;
	reg [0:0] injection_channels_173_;
	reg [0:0] injection_channels_172_;
	reg [0:0] injection_channels_171_;
	reg [0:0] injection_channels_170_;
	reg [0:0] injection_channels_169_;
	reg [0:0] injection_channels_168_;
	reg [0:0] injection_channels_167_;
	reg [0:0] injection_channels_166_;
	reg [0:0] injection_channels_165_;
	reg [0:0] injection_channels_164_;
	reg [0:0] injection_channels_163_;
	reg [0:0] injection_channels_162_;
	reg [0:0] injection_channels_161_;
	reg [0:0] injection_channels_160_;
	reg [0:0] injection_channels_159_;
	reg [0:0] injection_channels_158_;
	reg [0:0] injection_channels_157_;
	reg [0:0] injection_channels_156_;
	reg [0:0] injection_channels_155_;
	reg [0:0] injection_channels_154_;
	reg [0:0] injection_channels_153_;
	reg [0:0] injection_channels_152_;
	reg [0:0] injection_channels_151_;
	reg [0:0] injection_channels_150_;
	reg [0:0] injection_channels_149_;
	reg [0:0] injection_channels_148_;
	reg [0:0] injection_channels_147_;
	reg [0:0] injection_channels_146_;
	reg [0:0] injection_channels_145_;
	reg [0:0] injection_channels_144_;
	reg [0:0] injection_channels_143_;
	reg [0:0] injection_channels_142_;
	reg [0:0] injection_channels_141_;
	reg [0:0] injection_channels_140_;
	reg [0:0] injection_channels_139_;
	reg [0:0] injection_channels_138_;
	reg [0:0] injection_channels_137_;
	reg [0:0] injection_channels_136_;
	reg [0:0] injection_channels_135_;
	reg [0:0] injection_channels_134_;
	reg [0:0] injection_channels_133_;
	reg [0:0] injection_channels_132_;
	reg [0:0] injection_channels_131_;
	reg [0:0] injection_channels_130_;
	reg [0:0] injection_channels_129_;
	reg [0:0] injection_channels_128_;
	reg [0:0] injection_channels_127_;
	reg [0:0] injection_channels_126_;
	reg [0:0] injection_channels_125_;
	reg [0:0] injection_channels_124_;
	reg [0:0] injection_channels_123_;
	reg [0:0] injection_channels_122_;
	reg [0:0] injection_channels_121_;
	reg [0:0] injection_channels_120_;
	reg [0:0] injection_channels_119_;
	reg [0:0] injection_channels_118_;
	reg [0:0] injection_channels_117_;
	reg [0:0] injection_channels_116_;
	reg [0:0] injection_channels_115_;
	reg [0:0] injection_channels_114_;
	reg [0:0] injection_channels_113_;
	reg [0:0] injection_channels_112_;
	reg [0:0] injection_channels_111_;
	reg [0:0] injection_channels_110_;
	reg [0:0] injection_channels_109_;
	reg [0:0] injection_channels_108_;
	reg [0:0] injection_channels_107_;
	reg [0:0] injection_channels_106_;
	reg [0:0] injection_channels_105_;
	reg [0:0] injection_channels_104_;
	reg [0:0] injection_channels_103_;
	reg [0:0] injection_channels_102_;
	reg [0:0] injection_channels_101_;
	reg [0:0] injection_channels_100_;
	reg [0:0] injection_channels_99_;
	reg [0:0] injection_channels_98_;
	reg [0:0] injection_channels_97_;
	reg [0:0] injection_channels_96_;
	reg [0:0] injection_channels_95_;
	reg [0:0] injection_channels_94_;
	reg [0:0] injection_channels_93_;
	reg [0:0] injection_channels_92_;
	reg [0:0] injection_channels_91_;
	reg [0:0] injection_channels_90_;
	reg [0:0] injection_channels_89_;
	reg [0:0] injection_channels_88_;
	reg [0:0] injection_channels_87_;
	reg [0:0] injection_channels_86_;
	reg [0:0] injection_channels_85_;
	reg [0:0] injection_channels_84_;
	reg [0:0] injection_channels_83_;
	reg [0:0] injection_channels_82_;
	reg [0:0] injection_channels_81_;
	reg [0:0] injection_channels_80_;
	reg [0:0] injection_channels_79_;
	reg [0:0] injection_channels_78_;
	reg [0:0] injection_channels_77_;
	reg [0:0] injection_channels_76_;
	reg [0:0] injection_channels_75_;
	reg [0:0] injection_channels_74_;
	reg [0:0] injection_channels_73_;
	reg [0:0] injection_channels_72_;
	reg [0:0] injection_channels_71_;
	reg [0:0] injection_channels_70_;
	reg [0:0] injection_channels_69_;
	reg [0:0] injection_channels_68_;
	reg [0:0] injection_channels_67_;
	reg [0:0] injection_channels_66_;
	reg [0:0] injection_channels_65_;
	reg [0:0] injection_channels_64_;
	reg [0:0] injection_channels_63_;
	reg [0:0] injection_channels_62_;
	reg [0:0] injection_channels_61_;
	reg [0:0] injection_channels_60_;
	reg [0:0] injection_channels_59_;
	reg [0:0] injection_channels_58_;
	reg [0:0] injection_channels_57_;
	reg [0:0] injection_channels_56_;
	reg [0:0] injection_channels_55_;
	reg [0:0] injection_channels_54_;
	reg [0:0] injection_channels_53_;
	reg [0:0] injection_channels_52_;
	reg [0:0] injection_channels_51_;
	reg [0:0] injection_channels_50_;
	reg [0:0] injection_channels_49_;
	reg [0:0] injection_channels_48_;
	reg [0:0] injection_channels_47_;
	reg [0:0] injection_channels_46_;
	reg [0:0] injection_channels_45_;
	reg [0:0] injection_channels_44_;
	reg [0:0] injection_channels_43_;
	reg [0:0] injection_channels_42_;
	reg [0:0] injection_channels_41_;
	reg [0:0] injection_channels_40_;
	reg [0:0] injection_channels_39_;
	reg [0:0] injection_channels_38_;
	reg [0:0] injection_channels_37_;
	reg [0:0] injection_channels_36_;
	reg [0:0] injection_channels_35_;
	reg [0:0] injection_channels_34_;
	reg [0:0] injection_channels_33_;
	reg [0:0] injection_channels_32_;
	reg [0:0] injection_channels_31_;
	reg [0:0] injection_channels_30_;
	reg [0:0] injection_channels_29_;
	reg [0:0] injection_channels_28_;
	reg [0:0] injection_channels_27_;
	reg [0:0] injection_channels_26_;
	reg [0:0] injection_channels_25_;
	reg [0:0] injection_channels_24_;
	reg [0:0] injection_channels_23_;
	reg [0:0] injection_channels_22_;
	reg [0:0] injection_channels_21_;
	reg [0:0] injection_channels_20_;
	reg [0:0] injection_channels_19_;
	reg [0:0] injection_channels_18_;
	reg [0:0] injection_channels_17_;
	reg [0:0] injection_channels_16_;
	reg [0:0] injection_channels_15_;
	reg [0:0] injection_channels_14_;
	reg [0:0] injection_channels_13_;
	reg [0:0] injection_channels_12_;
	reg [0:0] injection_channels_11_;
	reg [0:0] injection_channels_10_;
	reg [0:0] injection_channels_9_;
	reg [0:0] injection_channels_8_;
	reg [0:0] injection_channels_7_;
	reg [0:0] injection_channels_6_;
	reg [0:0] injection_channels_5_;
	reg [0:0] injection_channels_4_;
	reg [0:0] injection_channels_3_;
	reg [0:0] injection_channels_2_;
	reg [0:0] injection_channels_1_;
	reg [0:0] injection_channels_0_;
	reg [0:0] ejection_flow_ctrl_26_;
	reg [0:0] ejection_flow_ctrl_25_;
	reg [0:0] ejection_flow_ctrl_24_;
	reg [0:0] ejection_flow_ctrl_23_;
	reg [0:0] ejection_flow_ctrl_22_;
	reg [0:0] ejection_flow_ctrl_21_;
	reg [0:0] ejection_flow_ctrl_20_;
	reg [0:0] ejection_flow_ctrl_19_;
	reg [0:0] ejection_flow_ctrl_18_;
	reg [0:0] ejection_flow_ctrl_17_;
	reg [0:0] ejection_flow_ctrl_16_;
	reg [0:0] ejection_flow_ctrl_15_;
	reg [0:0] ejection_flow_ctrl_14_;
	reg [0:0] ejection_flow_ctrl_13_;
	reg [0:0] ejection_flow_ctrl_12_;
	reg [0:0] ejection_flow_ctrl_11_;
	reg [0:0] ejection_flow_ctrl_10_;
	reg [0:0] ejection_flow_ctrl_9_;
	reg [0:0] ejection_flow_ctrl_8_;
	reg [0:0] ejection_flow_ctrl_7_;
	reg [0:0] ejection_flow_ctrl_6_;
	reg [0:0] ejection_flow_ctrl_5_;
	reg [0:0] ejection_flow_ctrl_4_;
	reg [0:0] ejection_flow_ctrl_3_;
	reg [0:0] ejection_flow_ctrl_2_;
	reg [0:0] ejection_flow_ctrl_1_;
	reg [0:0] ejection_flow_ctrl_0_;

// ----- FPGA fabric outputs -------
	wire [0:0] injection_flow_ctrl_26__gfpga;
	wire [0:0] injection_flow_ctrl_25__gfpga;
	wire [0:0] injection_flow_ctrl_24__gfpga;
	wire [0:0] injection_flow_ctrl_23__gfpga;
	wire [0:0] injection_flow_ctrl_22__gfpga;
	wire [0:0] injection_flow_ctrl_21__gfpga;
	wire [0:0] injection_flow_ctrl_20__gfpga;
	wire [0:0] injection_flow_ctrl_19__gfpga;
	wire [0:0] injection_flow_ctrl_18__gfpga;
	wire [0:0] injection_flow_ctrl_17__gfpga;
	wire [0:0] injection_flow_ctrl_16__gfpga;
	wire [0:0] injection_flow_ctrl_15__gfpga;
	wire [0:0] injection_flow_ctrl_14__gfpga;
	wire [0:0] injection_flow_ctrl_13__gfpga;
	wire [0:0] injection_flow_ctrl_12__gfpga;
	wire [0:0] injection_flow_ctrl_11__gfpga;
	wire [0:0] injection_flow_ctrl_10__gfpga;
	wire [0:0] injection_flow_ctrl_9__gfpga;
	wire [0:0] injection_flow_ctrl_8__gfpga;
	wire [0:0] injection_flow_ctrl_7__gfpga;
	wire [0:0] injection_flow_ctrl_6__gfpga;
	wire [0:0] injection_flow_ctrl_5__gfpga;
	wire [0:0] injection_flow_ctrl_4__gfpga;
	wire [0:0] injection_flow_ctrl_3__gfpga;
	wire [0:0] injection_flow_ctrl_2__gfpga;
	wire [0:0] injection_flow_ctrl_1__gfpga;
	wire [0:0] injection_flow_ctrl_0__gfpga;
	wire [0:0] ejection_channels_629__gfpga;
	wire [0:0] ejection_channels_628__gfpga;
	wire [0:0] ejection_channels_627__gfpga;
	wire [0:0] ejection_channels_626__gfpga;
	wire [0:0] ejection_channels_625__gfpga;
	wire [0:0] ejection_channels_624__gfpga;
	wire [0:0] ejection_channels_623__gfpga;
	wire [0:0] ejection_channels_622__gfpga;
	wire [0:0] ejection_channels_621__gfpga;
	wire [0:0] ejection_channels_620__gfpga;
	wire [0:0] ejection_channels_619__gfpga;
	wire [0:0] ejection_channels_618__gfpga;
	wire [0:0] ejection_channels_617__gfpga;
	wire [0:0] ejection_channels_616__gfpga;
	wire [0:0] ejection_channels_615__gfpga;
	wire [0:0] ejection_channels_614__gfpga;
	wire [0:0] ejection_channels_613__gfpga;
	wire [0:0] ejection_channels_612__gfpga;
	wire [0:0] ejection_channels_611__gfpga;
	wire [0:0] ejection_channels_610__gfpga;
	wire [0:0] ejection_channels_609__gfpga;
	wire [0:0] ejection_channels_608__gfpga;
	wire [0:0] ejection_channels_607__gfpga;
	wire [0:0] ejection_channels_606__gfpga;
	wire [0:0] ejection_channels_605__gfpga;
	wire [0:0] ejection_channels_604__gfpga;
	wire [0:0] ejection_channels_603__gfpga;
	wire [0:0] ejection_channels_602__gfpga;
	wire [0:0] ejection_channels_601__gfpga;
	wire [0:0] ejection_channels_600__gfpga;
	wire [0:0] ejection_channels_599__gfpga;
	wire [0:0] ejection_channels_598__gfpga;
	wire [0:0] ejection_channels_597__gfpga;
	wire [0:0] ejection_channels_596__gfpga;
	wire [0:0] ejection_channels_595__gfpga;
	wire [0:0] ejection_channels_594__gfpga;
	wire [0:0] ejection_channels_593__gfpga;
	wire [0:0] ejection_channels_592__gfpga;
	wire [0:0] ejection_channels_591__gfpga;
	wire [0:0] ejection_channels_590__gfpga;
	wire [0:0] ejection_channels_589__gfpga;
	wire [0:0] ejection_channels_588__gfpga;
	wire [0:0] ejection_channels_587__gfpga;
	wire [0:0] ejection_channels_586__gfpga;
	wire [0:0] ejection_channels_585__gfpga;
	wire [0:0] ejection_channels_584__gfpga;
	wire [0:0] ejection_channels_583__gfpga;
	wire [0:0] ejection_channels_582__gfpga;
	wire [0:0] ejection_channels_581__gfpga;
	wire [0:0] ejection_channels_580__gfpga;
	wire [0:0] ejection_channels_579__gfpga;
	wire [0:0] ejection_channels_578__gfpga;
	wire [0:0] ejection_channels_577__gfpga;
	wire [0:0] ejection_channels_576__gfpga;
	wire [0:0] ejection_channels_575__gfpga;
	wire [0:0] ejection_channels_574__gfpga;
	wire [0:0] ejection_channels_573__gfpga;
	wire [0:0] ejection_channels_572__gfpga;
	wire [0:0] ejection_channels_571__gfpga;
	wire [0:0] ejection_channels_570__gfpga;
	wire [0:0] ejection_channels_569__gfpga;
	wire [0:0] ejection_channels_568__gfpga;
	wire [0:0] ejection_channels_567__gfpga;
	wire [0:0] ejection_channels_566__gfpga;
	wire [0:0] ejection_channels_565__gfpga;
	wire [0:0] ejection_channels_564__gfpga;
	wire [0:0] ejection_channels_563__gfpga;
	wire [0:0] ejection_channels_562__gfpga;
	wire [0:0] ejection_channels_561__gfpga;
	wire [0:0] ejection_channels_560__gfpga;
	wire [0:0] ejection_channels_559__gfpga;
	wire [0:0] ejection_channels_558__gfpga;
	wire [0:0] ejection_channels_557__gfpga;
	wire [0:0] ejection_channels_556__gfpga;
	wire [0:0] ejection_channels_555__gfpga;
	wire [0:0] ejection_channels_554__gfpga;
	wire [0:0] ejection_channels_553__gfpga;
	wire [0:0] ejection_channels_552__gfpga;
	wire [0:0] ejection_channels_551__gfpga;
	wire [0:0] ejection_channels_550__gfpga;
	wire [0:0] ejection_channels_549__gfpga;
	wire [0:0] ejection_channels_548__gfpga;
	wire [0:0] ejection_channels_547__gfpga;
	wire [0:0] ejection_channels_546__gfpga;
	wire [0:0] ejection_channels_545__gfpga;
	wire [0:0] ejection_channels_544__gfpga;
	wire [0:0] ejection_channels_543__gfpga;
	wire [0:0] ejection_channels_542__gfpga;
	wire [0:0] ejection_channels_541__gfpga;
	wire [0:0] ejection_channels_540__gfpga;
	wire [0:0] ejection_channels_539__gfpga;
	wire [0:0] ejection_channels_538__gfpga;
	wire [0:0] ejection_channels_537__gfpga;
	wire [0:0] ejection_channels_536__gfpga;
	wire [0:0] ejection_channels_535__gfpga;
	wire [0:0] ejection_channels_534__gfpga;
	wire [0:0] ejection_channels_533__gfpga;
	wire [0:0] ejection_channels_532__gfpga;
	wire [0:0] ejection_channels_531__gfpga;
	wire [0:0] ejection_channels_530__gfpga;
	wire [0:0] ejection_channels_529__gfpga;
	wire [0:0] ejection_channels_528__gfpga;
	wire [0:0] ejection_channels_527__gfpga;
	wire [0:0] ejection_channels_526__gfpga;
	wire [0:0] ejection_channels_525__gfpga;
	wire [0:0] ejection_channels_524__gfpga;
	wire [0:0] ejection_channels_523__gfpga;
	wire [0:0] ejection_channels_522__gfpga;
	wire [0:0] ejection_channels_521__gfpga;
	wire [0:0] ejection_channels_520__gfpga;
	wire [0:0] ejection_channels_519__gfpga;
	wire [0:0] ejection_channels_518__gfpga;
	wire [0:0] ejection_channels_517__gfpga;
	wire [0:0] ejection_channels_516__gfpga;
	wire [0:0] ejection_channels_515__gfpga;
	wire [0:0] ejection_channels_514__gfpga;
	wire [0:0] ejection_channels_513__gfpga;
	wire [0:0] ejection_channels_512__gfpga;
	wire [0:0] ejection_channels_511__gfpga;
	wire [0:0] ejection_channels_510__gfpga;
	wire [0:0] ejection_channels_509__gfpga;
	wire [0:0] ejection_channels_508__gfpga;
	wire [0:0] ejection_channels_507__gfpga;
	wire [0:0] ejection_channels_506__gfpga;
	wire [0:0] ejection_channels_505__gfpga;
	wire [0:0] ejection_channels_504__gfpga;
	wire [0:0] ejection_channels_503__gfpga;
	wire [0:0] ejection_channels_502__gfpga;
	wire [0:0] ejection_channels_501__gfpga;
	wire [0:0] ejection_channels_500__gfpga;
	wire [0:0] ejection_channels_499__gfpga;
	wire [0:0] ejection_channels_498__gfpga;
	wire [0:0] ejection_channels_497__gfpga;
	wire [0:0] ejection_channels_496__gfpga;
	wire [0:0] ejection_channels_495__gfpga;
	wire [0:0] ejection_channels_494__gfpga;
	wire [0:0] ejection_channels_493__gfpga;
	wire [0:0] ejection_channels_492__gfpga;
	wire [0:0] ejection_channels_491__gfpga;
	wire [0:0] ejection_channels_490__gfpga;
	wire [0:0] ejection_channels_489__gfpga;
	wire [0:0] ejection_channels_488__gfpga;
	wire [0:0] ejection_channels_487__gfpga;
	wire [0:0] ejection_channels_486__gfpga;
	wire [0:0] ejection_channels_485__gfpga;
	wire [0:0] ejection_channels_484__gfpga;
	wire [0:0] ejection_channels_483__gfpga;
	wire [0:0] ejection_channels_482__gfpga;
	wire [0:0] ejection_channels_481__gfpga;
	wire [0:0] ejection_channels_480__gfpga;
	wire [0:0] ejection_channels_479__gfpga;
	wire [0:0] ejection_channels_478__gfpga;
	wire [0:0] ejection_channels_477__gfpga;
	wire [0:0] ejection_channels_476__gfpga;
	wire [0:0] ejection_channels_475__gfpga;
	wire [0:0] ejection_channels_474__gfpga;
	wire [0:0] ejection_channels_473__gfpga;
	wire [0:0] ejection_channels_472__gfpga;
	wire [0:0] ejection_channels_471__gfpga;
	wire [0:0] ejection_channels_470__gfpga;
	wire [0:0] ejection_channels_469__gfpga;
	wire [0:0] ejection_channels_468__gfpga;
	wire [0:0] ejection_channels_467__gfpga;
	wire [0:0] ejection_channels_466__gfpga;
	wire [0:0] ejection_channels_465__gfpga;
	wire [0:0] ejection_channels_464__gfpga;
	wire [0:0] ejection_channels_463__gfpga;
	wire [0:0] ejection_channels_462__gfpga;
	wire [0:0] ejection_channels_461__gfpga;
	wire [0:0] ejection_channels_460__gfpga;
	wire [0:0] ejection_channels_459__gfpga;
	wire [0:0] ejection_channels_458__gfpga;
	wire [0:0] ejection_channels_457__gfpga;
	wire [0:0] ejection_channels_456__gfpga;
	wire [0:0] ejection_channels_455__gfpga;
	wire [0:0] ejection_channels_454__gfpga;
	wire [0:0] ejection_channels_453__gfpga;
	wire [0:0] ejection_channels_452__gfpga;
	wire [0:0] ejection_channels_451__gfpga;
	wire [0:0] ejection_channels_450__gfpga;
	wire [0:0] ejection_channels_449__gfpga;
	wire [0:0] ejection_channels_448__gfpga;
	wire [0:0] ejection_channels_447__gfpga;
	wire [0:0] ejection_channels_446__gfpga;
	wire [0:0] ejection_channels_445__gfpga;
	wire [0:0] ejection_channels_444__gfpga;
	wire [0:0] ejection_channels_443__gfpga;
	wire [0:0] ejection_channels_442__gfpga;
	wire [0:0] ejection_channels_441__gfpga;
	wire [0:0] ejection_channels_440__gfpga;
	wire [0:0] ejection_channels_439__gfpga;
	wire [0:0] ejection_channels_438__gfpga;
	wire [0:0] ejection_channels_437__gfpga;
	wire [0:0] ejection_channels_436__gfpga;
	wire [0:0] ejection_channels_435__gfpga;
	wire [0:0] ejection_channels_434__gfpga;
	wire [0:0] ejection_channels_433__gfpga;
	wire [0:0] ejection_channels_432__gfpga;
	wire [0:0] ejection_channels_431__gfpga;
	wire [0:0] ejection_channels_430__gfpga;
	wire [0:0] ejection_channels_429__gfpga;
	wire [0:0] ejection_channels_428__gfpga;
	wire [0:0] ejection_channels_427__gfpga;
	wire [0:0] ejection_channels_426__gfpga;
	wire [0:0] ejection_channels_425__gfpga;
	wire [0:0] ejection_channels_424__gfpga;
	wire [0:0] ejection_channels_423__gfpga;
	wire [0:0] ejection_channels_422__gfpga;
	wire [0:0] ejection_channels_421__gfpga;
	wire [0:0] ejection_channels_420__gfpga;
	wire [0:0] ejection_channels_419__gfpga;
	wire [0:0] ejection_channels_418__gfpga;
	wire [0:0] ejection_channels_417__gfpga;
	wire [0:0] ejection_channels_416__gfpga;
	wire [0:0] ejection_channels_415__gfpga;
	wire [0:0] ejection_channels_414__gfpga;
	wire [0:0] ejection_channels_413__gfpga;
	wire [0:0] ejection_channels_412__gfpga;
	wire [0:0] ejection_channels_411__gfpga;
	wire [0:0] ejection_channels_410__gfpga;
	wire [0:0] ejection_channels_409__gfpga;
	wire [0:0] ejection_channels_408__gfpga;
	wire [0:0] ejection_channels_407__gfpga;
	wire [0:0] ejection_channels_406__gfpga;
	wire [0:0] ejection_channels_405__gfpga;
	wire [0:0] ejection_channels_404__gfpga;
	wire [0:0] ejection_channels_403__gfpga;
	wire [0:0] ejection_channels_402__gfpga;
	wire [0:0] ejection_channels_401__gfpga;
	wire [0:0] ejection_channels_400__gfpga;
	wire [0:0] ejection_channels_399__gfpga;
	wire [0:0] ejection_channels_398__gfpga;
	wire [0:0] ejection_channels_397__gfpga;
	wire [0:0] ejection_channels_396__gfpga;
	wire [0:0] ejection_channels_395__gfpga;
	wire [0:0] ejection_channels_394__gfpga;
	wire [0:0] ejection_channels_393__gfpga;
	wire [0:0] ejection_channels_392__gfpga;
	wire [0:0] ejection_channels_391__gfpga;
	wire [0:0] ejection_channels_390__gfpga;
	wire [0:0] ejection_channels_389__gfpga;
	wire [0:0] ejection_channels_388__gfpga;
	wire [0:0] ejection_channels_387__gfpga;
	wire [0:0] ejection_channels_386__gfpga;
	wire [0:0] ejection_channels_385__gfpga;
	wire [0:0] ejection_channels_384__gfpga;
	wire [0:0] ejection_channels_383__gfpga;
	wire [0:0] ejection_channels_382__gfpga;
	wire [0:0] ejection_channels_381__gfpga;
	wire [0:0] ejection_channels_380__gfpga;
	wire [0:0] ejection_channels_379__gfpga;
	wire [0:0] ejection_channels_378__gfpga;
	wire [0:0] ejection_channels_377__gfpga;
	wire [0:0] ejection_channels_376__gfpga;
	wire [0:0] ejection_channels_375__gfpga;
	wire [0:0] ejection_channels_374__gfpga;
	wire [0:0] ejection_channels_373__gfpga;
	wire [0:0] ejection_channels_372__gfpga;
	wire [0:0] ejection_channels_371__gfpga;
	wire [0:0] ejection_channels_370__gfpga;
	wire [0:0] ejection_channels_369__gfpga;
	wire [0:0] ejection_channels_368__gfpga;
	wire [0:0] ejection_channels_367__gfpga;
	wire [0:0] ejection_channels_366__gfpga;
	wire [0:0] ejection_channels_365__gfpga;
	wire [0:0] ejection_channels_364__gfpga;
	wire [0:0] ejection_channels_363__gfpga;
	wire [0:0] ejection_channels_362__gfpga;
	wire [0:0] ejection_channels_361__gfpga;
	wire [0:0] ejection_channels_360__gfpga;
	wire [0:0] ejection_channels_359__gfpga;
	wire [0:0] ejection_channels_358__gfpga;
	wire [0:0] ejection_channels_357__gfpga;
	wire [0:0] ejection_channels_356__gfpga;
	wire [0:0] ejection_channels_355__gfpga;
	wire [0:0] ejection_channels_354__gfpga;
	wire [0:0] ejection_channels_353__gfpga;
	wire [0:0] ejection_channels_352__gfpga;
	wire [0:0] ejection_channels_351__gfpga;
	wire [0:0] ejection_channels_350__gfpga;
	wire [0:0] ejection_channels_349__gfpga;
	wire [0:0] ejection_channels_348__gfpga;
	wire [0:0] ejection_channels_347__gfpga;
	wire [0:0] ejection_channels_346__gfpga;
	wire [0:0] ejection_channels_345__gfpga;
	wire [0:0] ejection_channels_344__gfpga;
	wire [0:0] ejection_channels_343__gfpga;
	wire [0:0] ejection_channels_342__gfpga;
	wire [0:0] ejection_channels_341__gfpga;
	wire [0:0] ejection_channels_340__gfpga;
	wire [0:0] ejection_channels_339__gfpga;
	wire [0:0] ejection_channels_338__gfpga;
	wire [0:0] ejection_channels_337__gfpga;
	wire [0:0] ejection_channels_336__gfpga;
	wire [0:0] ejection_channels_335__gfpga;
	wire [0:0] ejection_channels_334__gfpga;
	wire [0:0] ejection_channels_333__gfpga;
	wire [0:0] ejection_channels_332__gfpga;
	wire [0:0] ejection_channels_331__gfpga;
	wire [0:0] ejection_channels_330__gfpga;
	wire [0:0] ejection_channels_329__gfpga;
	wire [0:0] ejection_channels_328__gfpga;
	wire [0:0] ejection_channels_327__gfpga;
	wire [0:0] ejection_channels_326__gfpga;
	wire [0:0] ejection_channels_325__gfpga;
	wire [0:0] ejection_channels_324__gfpga;
	wire [0:0] ejection_channels_323__gfpga;
	wire [0:0] ejection_channels_322__gfpga;
	wire [0:0] ejection_channels_321__gfpga;
	wire [0:0] ejection_channels_320__gfpga;
	wire [0:0] ejection_channels_319__gfpga;
	wire [0:0] ejection_channels_318__gfpga;
	wire [0:0] ejection_channels_317__gfpga;
	wire [0:0] ejection_channels_316__gfpga;
	wire [0:0] ejection_channels_315__gfpga;
	wire [0:0] ejection_channels_314__gfpga;
	wire [0:0] ejection_channels_313__gfpga;
	wire [0:0] ejection_channels_312__gfpga;
	wire [0:0] ejection_channels_311__gfpga;
	wire [0:0] ejection_channels_310__gfpga;
	wire [0:0] ejection_channels_309__gfpga;
	wire [0:0] ejection_channels_308__gfpga;
	wire [0:0] ejection_channels_307__gfpga;
	wire [0:0] ejection_channels_306__gfpga;
	wire [0:0] ejection_channels_305__gfpga;
	wire [0:0] ejection_channels_304__gfpga;
	wire [0:0] ejection_channels_303__gfpga;
	wire [0:0] ejection_channels_302__gfpga;
	wire [0:0] ejection_channels_301__gfpga;
	wire [0:0] ejection_channels_300__gfpga;
	wire [0:0] ejection_channels_299__gfpga;
	wire [0:0] ejection_channels_298__gfpga;
	wire [0:0] ejection_channels_297__gfpga;
	wire [0:0] ejection_channels_296__gfpga;
	wire [0:0] ejection_channels_295__gfpga;
	wire [0:0] ejection_channels_294__gfpga;
	wire [0:0] ejection_channels_293__gfpga;
	wire [0:0] ejection_channels_292__gfpga;
	wire [0:0] ejection_channels_291__gfpga;
	wire [0:0] ejection_channels_290__gfpga;
	wire [0:0] ejection_channels_289__gfpga;
	wire [0:0] ejection_channels_288__gfpga;
	wire [0:0] ejection_channels_287__gfpga;
	wire [0:0] ejection_channels_286__gfpga;
	wire [0:0] ejection_channels_285__gfpga;
	wire [0:0] ejection_channels_284__gfpga;
	wire [0:0] ejection_channels_283__gfpga;
	wire [0:0] ejection_channels_282__gfpga;
	wire [0:0] ejection_channels_281__gfpga;
	wire [0:0] ejection_channels_280__gfpga;
	wire [0:0] ejection_channels_279__gfpga;
	wire [0:0] ejection_channels_278__gfpga;
	wire [0:0] ejection_channels_277__gfpga;
	wire [0:0] ejection_channels_276__gfpga;
	wire [0:0] ejection_channels_275__gfpga;
	wire [0:0] ejection_channels_274__gfpga;
	wire [0:0] ejection_channels_273__gfpga;
	wire [0:0] ejection_channels_272__gfpga;
	wire [0:0] ejection_channels_271__gfpga;
	wire [0:0] ejection_channels_270__gfpga;
	wire [0:0] ejection_channels_269__gfpga;
	wire [0:0] ejection_channels_268__gfpga;
	wire [0:0] ejection_channels_267__gfpga;
	wire [0:0] ejection_channels_266__gfpga;
	wire [0:0] ejection_channels_265__gfpga;
	wire [0:0] ejection_channels_264__gfpga;
	wire [0:0] ejection_channels_263__gfpga;
	wire [0:0] ejection_channels_262__gfpga;
	wire [0:0] ejection_channels_261__gfpga;
	wire [0:0] ejection_channels_260__gfpga;
	wire [0:0] ejection_channels_259__gfpga;
	wire [0:0] ejection_channels_258__gfpga;
	wire [0:0] ejection_channels_257__gfpga;
	wire [0:0] ejection_channels_256__gfpga;
	wire [0:0] ejection_channels_255__gfpga;
	wire [0:0] ejection_channels_254__gfpga;
	wire [0:0] ejection_channels_253__gfpga;
	wire [0:0] ejection_channels_252__gfpga;
	wire [0:0] ejection_channels_251__gfpga;
	wire [0:0] ejection_channels_250__gfpga;
	wire [0:0] ejection_channels_249__gfpga;
	wire [0:0] ejection_channels_248__gfpga;
	wire [0:0] ejection_channels_247__gfpga;
	wire [0:0] ejection_channels_246__gfpga;
	wire [0:0] ejection_channels_245__gfpga;
	wire [0:0] ejection_channels_244__gfpga;
	wire [0:0] ejection_channels_243__gfpga;
	wire [0:0] ejection_channels_242__gfpga;
	wire [0:0] ejection_channels_241__gfpga;
	wire [0:0] ejection_channels_240__gfpga;
	wire [0:0] ejection_channels_239__gfpga;
	wire [0:0] ejection_channels_238__gfpga;
	wire [0:0] ejection_channels_237__gfpga;
	wire [0:0] ejection_channels_236__gfpga;
	wire [0:0] ejection_channels_235__gfpga;
	wire [0:0] ejection_channels_234__gfpga;
	wire [0:0] ejection_channels_233__gfpga;
	wire [0:0] ejection_channels_232__gfpga;
	wire [0:0] ejection_channels_231__gfpga;
	wire [0:0] ejection_channels_230__gfpga;
	wire [0:0] ejection_channels_229__gfpga;
	wire [0:0] ejection_channels_228__gfpga;
	wire [0:0] ejection_channels_227__gfpga;
	wire [0:0] ejection_channels_226__gfpga;
	wire [0:0] ejection_channels_225__gfpga;
	wire [0:0] ejection_channels_224__gfpga;
	wire [0:0] ejection_channels_223__gfpga;
	wire [0:0] ejection_channels_222__gfpga;
	wire [0:0] ejection_channels_221__gfpga;
	wire [0:0] ejection_channels_220__gfpga;
	wire [0:0] ejection_channels_219__gfpga;
	wire [0:0] ejection_channels_218__gfpga;
	wire [0:0] ejection_channels_217__gfpga;
	wire [0:0] ejection_channels_216__gfpga;
	wire [0:0] ejection_channels_215__gfpga;
	wire [0:0] ejection_channels_214__gfpga;
	wire [0:0] ejection_channels_213__gfpga;
	wire [0:0] ejection_channels_212__gfpga;
	wire [0:0] ejection_channels_211__gfpga;
	wire [0:0] ejection_channels_210__gfpga;
	wire [0:0] ejection_channels_209__gfpga;
	wire [0:0] ejection_channels_208__gfpga;
	wire [0:0] ejection_channels_207__gfpga;
	wire [0:0] ejection_channels_206__gfpga;
	wire [0:0] ejection_channels_205__gfpga;
	wire [0:0] ejection_channels_204__gfpga;
	wire [0:0] ejection_channels_203__gfpga;
	wire [0:0] ejection_channels_202__gfpga;
	wire [0:0] ejection_channels_201__gfpga;
	wire [0:0] ejection_channels_200__gfpga;
	wire [0:0] ejection_channels_199__gfpga;
	wire [0:0] ejection_channels_198__gfpga;
	wire [0:0] ejection_channels_197__gfpga;
	wire [0:0] ejection_channels_196__gfpga;
	wire [0:0] ejection_channels_195__gfpga;
	wire [0:0] ejection_channels_194__gfpga;
	wire [0:0] ejection_channels_193__gfpga;
	wire [0:0] ejection_channels_192__gfpga;
	wire [0:0] ejection_channels_191__gfpga;
	wire [0:0] ejection_channels_190__gfpga;
	wire [0:0] ejection_channels_189__gfpga;
	wire [0:0] ejection_channels_188__gfpga;
	wire [0:0] ejection_channels_187__gfpga;
	wire [0:0] ejection_channels_186__gfpga;
	wire [0:0] ejection_channels_185__gfpga;
	wire [0:0] ejection_channels_184__gfpga;
	wire [0:0] ejection_channels_183__gfpga;
	wire [0:0] ejection_channels_182__gfpga;
	wire [0:0] ejection_channels_181__gfpga;
	wire [0:0] ejection_channels_180__gfpga;
	wire [0:0] ejection_channels_179__gfpga;
	wire [0:0] ejection_channels_178__gfpga;
	wire [0:0] ejection_channels_177__gfpga;
	wire [0:0] ejection_channels_176__gfpga;
	wire [0:0] ejection_channels_175__gfpga;
	wire [0:0] ejection_channels_174__gfpga;
	wire [0:0] ejection_channels_173__gfpga;
	wire [0:0] ejection_channels_172__gfpga;
	wire [0:0] ejection_channels_171__gfpga;
	wire [0:0] ejection_channels_170__gfpga;
	wire [0:0] ejection_channels_169__gfpga;
	wire [0:0] ejection_channels_168__gfpga;
	wire [0:0] ejection_channels_167__gfpga;
	wire [0:0] ejection_channels_166__gfpga;
	wire [0:0] ejection_channels_165__gfpga;
	wire [0:0] ejection_channels_164__gfpga;
	wire [0:0] ejection_channels_163__gfpga;
	wire [0:0] ejection_channels_162__gfpga;
	wire [0:0] ejection_channels_161__gfpga;
	wire [0:0] ejection_channels_160__gfpga;
	wire [0:0] ejection_channels_159__gfpga;
	wire [0:0] ejection_channels_158__gfpga;
	wire [0:0] ejection_channels_157__gfpga;
	wire [0:0] ejection_channels_156__gfpga;
	wire [0:0] ejection_channels_155__gfpga;
	wire [0:0] ejection_channels_154__gfpga;
	wire [0:0] ejection_channels_153__gfpga;
	wire [0:0] ejection_channels_152__gfpga;
	wire [0:0] ejection_channels_151__gfpga;
	wire [0:0] ejection_channels_150__gfpga;
	wire [0:0] ejection_channels_149__gfpga;
	wire [0:0] ejection_channels_148__gfpga;
	wire [0:0] ejection_channels_147__gfpga;
	wire [0:0] ejection_channels_146__gfpga;
	wire [0:0] ejection_channels_145__gfpga;
	wire [0:0] ejection_channels_144__gfpga;
	wire [0:0] ejection_channels_143__gfpga;
	wire [0:0] ejection_channels_142__gfpga;
	wire [0:0] ejection_channels_141__gfpga;
	wire [0:0] ejection_channels_140__gfpga;
	wire [0:0] ejection_channels_139__gfpga;
	wire [0:0] ejection_channels_138__gfpga;
	wire [0:0] ejection_channels_137__gfpga;
	wire [0:0] ejection_channels_136__gfpga;
	wire [0:0] ejection_channels_135__gfpga;
	wire [0:0] ejection_channels_134__gfpga;
	wire [0:0] ejection_channels_133__gfpga;
	wire [0:0] ejection_channels_132__gfpga;
	wire [0:0] ejection_channels_131__gfpga;
	wire [0:0] ejection_channels_130__gfpga;
	wire [0:0] ejection_channels_129__gfpga;
	wire [0:0] ejection_channels_128__gfpga;
	wire [0:0] ejection_channels_127__gfpga;
	wire [0:0] ejection_channels_126__gfpga;
	wire [0:0] ejection_channels_125__gfpga;
	wire [0:0] ejection_channels_124__gfpga;
	wire [0:0] ejection_channels_123__gfpga;
	wire [0:0] ejection_channels_122__gfpga;
	wire [0:0] ejection_channels_121__gfpga;
	wire [0:0] ejection_channels_120__gfpga;
	wire [0:0] ejection_channels_119__gfpga;
	wire [0:0] ejection_channels_118__gfpga;
	wire [0:0] ejection_channels_117__gfpga;
	wire [0:0] ejection_channels_116__gfpga;
	wire [0:0] ejection_channels_115__gfpga;
	wire [0:0] ejection_channels_114__gfpga;
	wire [0:0] ejection_channels_113__gfpga;
	wire [0:0] ejection_channels_112__gfpga;
	wire [0:0] ejection_channels_111__gfpga;
	wire [0:0] ejection_channels_110__gfpga;
	wire [0:0] ejection_channels_109__gfpga;
	wire [0:0] ejection_channels_108__gfpga;
	wire [0:0] ejection_channels_107__gfpga;
	wire [0:0] ejection_channels_106__gfpga;
	wire [0:0] ejection_channels_105__gfpga;
	wire [0:0] ejection_channels_104__gfpga;
	wire [0:0] ejection_channels_103__gfpga;
	wire [0:0] ejection_channels_102__gfpga;
	wire [0:0] ejection_channels_101__gfpga;
	wire [0:0] ejection_channels_100__gfpga;
	wire [0:0] ejection_channels_99__gfpga;
	wire [0:0] ejection_channels_98__gfpga;
	wire [0:0] ejection_channels_97__gfpga;
	wire [0:0] ejection_channels_96__gfpga;
	wire [0:0] ejection_channels_95__gfpga;
	wire [0:0] ejection_channels_94__gfpga;
	wire [0:0] ejection_channels_93__gfpga;
	wire [0:0] ejection_channels_92__gfpga;
	wire [0:0] ejection_channels_91__gfpga;
	wire [0:0] ejection_channels_90__gfpga;
	wire [0:0] ejection_channels_89__gfpga;
	wire [0:0] ejection_channels_88__gfpga;
	wire [0:0] ejection_channels_87__gfpga;
	wire [0:0] ejection_channels_86__gfpga;
	wire [0:0] ejection_channels_85__gfpga;
	wire [0:0] ejection_channels_84__gfpga;
	wire [0:0] ejection_channels_83__gfpga;
	wire [0:0] ejection_channels_82__gfpga;
	wire [0:0] ejection_channels_81__gfpga;
	wire [0:0] ejection_channels_80__gfpga;
	wire [0:0] ejection_channels_79__gfpga;
	wire [0:0] ejection_channels_78__gfpga;
	wire [0:0] ejection_channels_77__gfpga;
	wire [0:0] ejection_channels_76__gfpga;
	wire [0:0] ejection_channels_75__gfpga;
	wire [0:0] ejection_channels_74__gfpga;
	wire [0:0] ejection_channels_73__gfpga;
	wire [0:0] ejection_channels_72__gfpga;
	wire [0:0] ejection_channels_71__gfpga;
	wire [0:0] ejection_channels_70__gfpga;
	wire [0:0] ejection_channels_69__gfpga;
	wire [0:0] ejection_channels_68__gfpga;
	wire [0:0] ejection_channels_67__gfpga;
	wire [0:0] ejection_channels_66__gfpga;
	wire [0:0] ejection_channels_65__gfpga;
	wire [0:0] ejection_channels_64__gfpga;
	wire [0:0] ejection_channels_63__gfpga;
	wire [0:0] ejection_channels_62__gfpga;
	wire [0:0] ejection_channels_61__gfpga;
	wire [0:0] ejection_channels_60__gfpga;
	wire [0:0] ejection_channels_59__gfpga;
	wire [0:0] ejection_channels_58__gfpga;
	wire [0:0] ejection_channels_57__gfpga;
	wire [0:0] ejection_channels_56__gfpga;
	wire [0:0] ejection_channels_55__gfpga;
	wire [0:0] ejection_channels_54__gfpga;
	wire [0:0] ejection_channels_53__gfpga;
	wire [0:0] ejection_channels_52__gfpga;
	wire [0:0] ejection_channels_51__gfpga;
	wire [0:0] ejection_channels_50__gfpga;
	wire [0:0] ejection_channels_49__gfpga;
	wire [0:0] ejection_channels_48__gfpga;
	wire [0:0] ejection_channels_47__gfpga;
	wire [0:0] ejection_channels_46__gfpga;
	wire [0:0] ejection_channels_45__gfpga;
	wire [0:0] ejection_channels_44__gfpga;
	wire [0:0] ejection_channels_43__gfpga;
	wire [0:0] ejection_channels_42__gfpga;
	wire [0:0] ejection_channels_41__gfpga;
	wire [0:0] ejection_channels_40__gfpga;
	wire [0:0] ejection_channels_39__gfpga;
	wire [0:0] ejection_channels_38__gfpga;
	wire [0:0] ejection_channels_37__gfpga;
	wire [0:0] ejection_channels_36__gfpga;
	wire [0:0] ejection_channels_35__gfpga;
	wire [0:0] ejection_channels_34__gfpga;
	wire [0:0] ejection_channels_33__gfpga;
	wire [0:0] ejection_channels_32__gfpga;
	wire [0:0] ejection_channels_31__gfpga;
	wire [0:0] ejection_channels_30__gfpga;
	wire [0:0] ejection_channels_29__gfpga;
	wire [0:0] ejection_channels_28__gfpga;
	wire [0:0] ejection_channels_27__gfpga;
	wire [0:0] ejection_channels_26__gfpga;
	wire [0:0] ejection_channels_25__gfpga;
	wire [0:0] ejection_channels_24__gfpga;
	wire [0:0] ejection_channels_23__gfpga;
	wire [0:0] ejection_channels_22__gfpga;
	wire [0:0] ejection_channels_21__gfpga;
	wire [0:0] ejection_channels_20__gfpga;
	wire [0:0] ejection_channels_19__gfpga;
	wire [0:0] ejection_channels_18__gfpga;
	wire [0:0] ejection_channels_17__gfpga;
	wire [0:0] ejection_channels_16__gfpga;
	wire [0:0] ejection_channels_15__gfpga;
	wire [0:0] ejection_channels_14__gfpga;
	wire [0:0] ejection_channels_13__gfpga;
	wire [0:0] ejection_channels_12__gfpga;
	wire [0:0] ejection_channels_11__gfpga;
	wire [0:0] ejection_channels_10__gfpga;
	wire [0:0] ejection_channels_9__gfpga;
	wire [0:0] ejection_channels_8__gfpga;
	wire [0:0] ejection_channels_7__gfpga;
	wire [0:0] ejection_channels_6__gfpga;
	wire [0:0] ejection_channels_5__gfpga;
	wire [0:0] ejection_channels_4__gfpga;
	wire [0:0] ejection_channels_3__gfpga;
	wire [0:0] ejection_channels_2__gfpga;
	wire [0:0] ejection_channels_1__gfpga;
	wire [0:0] ejection_channels_0__gfpga;
	wire [0:0] rtr_error_8__gfpga;
	wire [0:0] rtr_error_7__gfpga;
	wire [0:0] rtr_error_6__gfpga;
	wire [0:0] rtr_error_5__gfpga;
	wire [0:0] rtr_error_4__gfpga;
	wire [0:0] rtr_error_3__gfpga;
	wire [0:0] rtr_error_2__gfpga;
	wire [0:0] rtr_error_1__gfpga;
	wire [0:0] rtr_error_0__gfpga;

// ----- Benchmark outputs -------
	wire [0:0] injection_flow_ctrl_26__bench;
	wire [0:0] injection_flow_ctrl_25__bench;
	wire [0:0] injection_flow_ctrl_24__bench;
	wire [0:0] injection_flow_ctrl_23__bench;
	wire [0:0] injection_flow_ctrl_22__bench;
	wire [0:0] injection_flow_ctrl_21__bench;
	wire [0:0] injection_flow_ctrl_20__bench;
	wire [0:0] injection_flow_ctrl_19__bench;
	wire [0:0] injection_flow_ctrl_18__bench;
	wire [0:0] injection_flow_ctrl_17__bench;
	wire [0:0] injection_flow_ctrl_16__bench;
	wire [0:0] injection_flow_ctrl_15__bench;
	wire [0:0] injection_flow_ctrl_14__bench;
	wire [0:0] injection_flow_ctrl_13__bench;
	wire [0:0] injection_flow_ctrl_12__bench;
	wire [0:0] injection_flow_ctrl_11__bench;
	wire [0:0] injection_flow_ctrl_10__bench;
	wire [0:0] injection_flow_ctrl_9__bench;
	wire [0:0] injection_flow_ctrl_8__bench;
	wire [0:0] injection_flow_ctrl_7__bench;
	wire [0:0] injection_flow_ctrl_6__bench;
	wire [0:0] injection_flow_ctrl_5__bench;
	wire [0:0] injection_flow_ctrl_4__bench;
	wire [0:0] injection_flow_ctrl_3__bench;
	wire [0:0] injection_flow_ctrl_2__bench;
	wire [0:0] injection_flow_ctrl_1__bench;
	wire [0:0] injection_flow_ctrl_0__bench;
	wire [0:0] ejection_channels_629__bench;
	wire [0:0] ejection_channels_628__bench;
	wire [0:0] ejection_channels_627__bench;
	wire [0:0] ejection_channels_626__bench;
	wire [0:0] ejection_channels_625__bench;
	wire [0:0] ejection_channels_624__bench;
	wire [0:0] ejection_channels_623__bench;
	wire [0:0] ejection_channels_622__bench;
	wire [0:0] ejection_channels_621__bench;
	wire [0:0] ejection_channels_620__bench;
	wire [0:0] ejection_channels_619__bench;
	wire [0:0] ejection_channels_618__bench;
	wire [0:0] ejection_channels_617__bench;
	wire [0:0] ejection_channels_616__bench;
	wire [0:0] ejection_channels_615__bench;
	wire [0:0] ejection_channels_614__bench;
	wire [0:0] ejection_channels_613__bench;
	wire [0:0] ejection_channels_612__bench;
	wire [0:0] ejection_channels_611__bench;
	wire [0:0] ejection_channels_610__bench;
	wire [0:0] ejection_channels_609__bench;
	wire [0:0] ejection_channels_608__bench;
	wire [0:0] ejection_channels_607__bench;
	wire [0:0] ejection_channels_606__bench;
	wire [0:0] ejection_channels_605__bench;
	wire [0:0] ejection_channels_604__bench;
	wire [0:0] ejection_channels_603__bench;
	wire [0:0] ejection_channels_602__bench;
	wire [0:0] ejection_channels_601__bench;
	wire [0:0] ejection_channels_600__bench;
	wire [0:0] ejection_channels_599__bench;
	wire [0:0] ejection_channels_598__bench;
	wire [0:0] ejection_channels_597__bench;
	wire [0:0] ejection_channels_596__bench;
	wire [0:0] ejection_channels_595__bench;
	wire [0:0] ejection_channels_594__bench;
	wire [0:0] ejection_channels_593__bench;
	wire [0:0] ejection_channels_592__bench;
	wire [0:0] ejection_channels_591__bench;
	wire [0:0] ejection_channels_590__bench;
	wire [0:0] ejection_channels_589__bench;
	wire [0:0] ejection_channels_588__bench;
	wire [0:0] ejection_channels_587__bench;
	wire [0:0] ejection_channels_586__bench;
	wire [0:0] ejection_channels_585__bench;
	wire [0:0] ejection_channels_584__bench;
	wire [0:0] ejection_channels_583__bench;
	wire [0:0] ejection_channels_582__bench;
	wire [0:0] ejection_channels_581__bench;
	wire [0:0] ejection_channels_580__bench;
	wire [0:0] ejection_channels_579__bench;
	wire [0:0] ejection_channels_578__bench;
	wire [0:0] ejection_channels_577__bench;
	wire [0:0] ejection_channels_576__bench;
	wire [0:0] ejection_channels_575__bench;
	wire [0:0] ejection_channels_574__bench;
	wire [0:0] ejection_channels_573__bench;
	wire [0:0] ejection_channels_572__bench;
	wire [0:0] ejection_channels_571__bench;
	wire [0:0] ejection_channels_570__bench;
	wire [0:0] ejection_channels_569__bench;
	wire [0:0] ejection_channels_568__bench;
	wire [0:0] ejection_channels_567__bench;
	wire [0:0] ejection_channels_566__bench;
	wire [0:0] ejection_channels_565__bench;
	wire [0:0] ejection_channels_564__bench;
	wire [0:0] ejection_channels_563__bench;
	wire [0:0] ejection_channels_562__bench;
	wire [0:0] ejection_channels_561__bench;
	wire [0:0] ejection_channels_560__bench;
	wire [0:0] ejection_channels_559__bench;
	wire [0:0] ejection_channels_558__bench;
	wire [0:0] ejection_channels_557__bench;
	wire [0:0] ejection_channels_556__bench;
	wire [0:0] ejection_channels_555__bench;
	wire [0:0] ejection_channels_554__bench;
	wire [0:0] ejection_channels_553__bench;
	wire [0:0] ejection_channels_552__bench;
	wire [0:0] ejection_channels_551__bench;
	wire [0:0] ejection_channels_550__bench;
	wire [0:0] ejection_channels_549__bench;
	wire [0:0] ejection_channels_548__bench;
	wire [0:0] ejection_channels_547__bench;
	wire [0:0] ejection_channels_546__bench;
	wire [0:0] ejection_channels_545__bench;
	wire [0:0] ejection_channels_544__bench;
	wire [0:0] ejection_channels_543__bench;
	wire [0:0] ejection_channels_542__bench;
	wire [0:0] ejection_channels_541__bench;
	wire [0:0] ejection_channels_540__bench;
	wire [0:0] ejection_channels_539__bench;
	wire [0:0] ejection_channels_538__bench;
	wire [0:0] ejection_channels_537__bench;
	wire [0:0] ejection_channels_536__bench;
	wire [0:0] ejection_channels_535__bench;
	wire [0:0] ejection_channels_534__bench;
	wire [0:0] ejection_channels_533__bench;
	wire [0:0] ejection_channels_532__bench;
	wire [0:0] ejection_channels_531__bench;
	wire [0:0] ejection_channels_530__bench;
	wire [0:0] ejection_channels_529__bench;
	wire [0:0] ejection_channels_528__bench;
	wire [0:0] ejection_channels_527__bench;
	wire [0:0] ejection_channels_526__bench;
	wire [0:0] ejection_channels_525__bench;
	wire [0:0] ejection_channels_524__bench;
	wire [0:0] ejection_channels_523__bench;
	wire [0:0] ejection_channels_522__bench;
	wire [0:0] ejection_channels_521__bench;
	wire [0:0] ejection_channels_520__bench;
	wire [0:0] ejection_channels_519__bench;
	wire [0:0] ejection_channels_518__bench;
	wire [0:0] ejection_channels_517__bench;
	wire [0:0] ejection_channels_516__bench;
	wire [0:0] ejection_channels_515__bench;
	wire [0:0] ejection_channels_514__bench;
	wire [0:0] ejection_channels_513__bench;
	wire [0:0] ejection_channels_512__bench;
	wire [0:0] ejection_channels_511__bench;
	wire [0:0] ejection_channels_510__bench;
	wire [0:0] ejection_channels_509__bench;
	wire [0:0] ejection_channels_508__bench;
	wire [0:0] ejection_channels_507__bench;
	wire [0:0] ejection_channels_506__bench;
	wire [0:0] ejection_channels_505__bench;
	wire [0:0] ejection_channels_504__bench;
	wire [0:0] ejection_channels_503__bench;
	wire [0:0] ejection_channels_502__bench;
	wire [0:0] ejection_channels_501__bench;
	wire [0:0] ejection_channels_500__bench;
	wire [0:0] ejection_channels_499__bench;
	wire [0:0] ejection_channels_498__bench;
	wire [0:0] ejection_channels_497__bench;
	wire [0:0] ejection_channels_496__bench;
	wire [0:0] ejection_channels_495__bench;
	wire [0:0] ejection_channels_494__bench;
	wire [0:0] ejection_channels_493__bench;
	wire [0:0] ejection_channels_492__bench;
	wire [0:0] ejection_channels_491__bench;
	wire [0:0] ejection_channels_490__bench;
	wire [0:0] ejection_channels_489__bench;
	wire [0:0] ejection_channels_488__bench;
	wire [0:0] ejection_channels_487__bench;
	wire [0:0] ejection_channels_486__bench;
	wire [0:0] ejection_channels_485__bench;
	wire [0:0] ejection_channels_484__bench;
	wire [0:0] ejection_channels_483__bench;
	wire [0:0] ejection_channels_482__bench;
	wire [0:0] ejection_channels_481__bench;
	wire [0:0] ejection_channels_480__bench;
	wire [0:0] ejection_channels_479__bench;
	wire [0:0] ejection_channels_478__bench;
	wire [0:0] ejection_channels_477__bench;
	wire [0:0] ejection_channels_476__bench;
	wire [0:0] ejection_channels_475__bench;
	wire [0:0] ejection_channels_474__bench;
	wire [0:0] ejection_channels_473__bench;
	wire [0:0] ejection_channels_472__bench;
	wire [0:0] ejection_channels_471__bench;
	wire [0:0] ejection_channels_470__bench;
	wire [0:0] ejection_channels_469__bench;
	wire [0:0] ejection_channels_468__bench;
	wire [0:0] ejection_channels_467__bench;
	wire [0:0] ejection_channels_466__bench;
	wire [0:0] ejection_channels_465__bench;
	wire [0:0] ejection_channels_464__bench;
	wire [0:0] ejection_channels_463__bench;
	wire [0:0] ejection_channels_462__bench;
	wire [0:0] ejection_channels_461__bench;
	wire [0:0] ejection_channels_460__bench;
	wire [0:0] ejection_channels_459__bench;
	wire [0:0] ejection_channels_458__bench;
	wire [0:0] ejection_channels_457__bench;
	wire [0:0] ejection_channels_456__bench;
	wire [0:0] ejection_channels_455__bench;
	wire [0:0] ejection_channels_454__bench;
	wire [0:0] ejection_channels_453__bench;
	wire [0:0] ejection_channels_452__bench;
	wire [0:0] ejection_channels_451__bench;
	wire [0:0] ejection_channels_450__bench;
	wire [0:0] ejection_channels_449__bench;
	wire [0:0] ejection_channels_448__bench;
	wire [0:0] ejection_channels_447__bench;
	wire [0:0] ejection_channels_446__bench;
	wire [0:0] ejection_channels_445__bench;
	wire [0:0] ejection_channels_444__bench;
	wire [0:0] ejection_channels_443__bench;
	wire [0:0] ejection_channels_442__bench;
	wire [0:0] ejection_channels_441__bench;
	wire [0:0] ejection_channels_440__bench;
	wire [0:0] ejection_channels_439__bench;
	wire [0:0] ejection_channels_438__bench;
	wire [0:0] ejection_channels_437__bench;
	wire [0:0] ejection_channels_436__bench;
	wire [0:0] ejection_channels_435__bench;
	wire [0:0] ejection_channels_434__bench;
	wire [0:0] ejection_channels_433__bench;
	wire [0:0] ejection_channels_432__bench;
	wire [0:0] ejection_channels_431__bench;
	wire [0:0] ejection_channels_430__bench;
	wire [0:0] ejection_channels_429__bench;
	wire [0:0] ejection_channels_428__bench;
	wire [0:0] ejection_channels_427__bench;
	wire [0:0] ejection_channels_426__bench;
	wire [0:0] ejection_channels_425__bench;
	wire [0:0] ejection_channels_424__bench;
	wire [0:0] ejection_channels_423__bench;
	wire [0:0] ejection_channels_422__bench;
	wire [0:0] ejection_channels_421__bench;
	wire [0:0] ejection_channels_420__bench;
	wire [0:0] ejection_channels_419__bench;
	wire [0:0] ejection_channels_418__bench;
	wire [0:0] ejection_channels_417__bench;
	wire [0:0] ejection_channels_416__bench;
	wire [0:0] ejection_channels_415__bench;
	wire [0:0] ejection_channels_414__bench;
	wire [0:0] ejection_channels_413__bench;
	wire [0:0] ejection_channels_412__bench;
	wire [0:0] ejection_channels_411__bench;
	wire [0:0] ejection_channels_410__bench;
	wire [0:0] ejection_channels_409__bench;
	wire [0:0] ejection_channels_408__bench;
	wire [0:0] ejection_channels_407__bench;
	wire [0:0] ejection_channels_406__bench;
	wire [0:0] ejection_channels_405__bench;
	wire [0:0] ejection_channels_404__bench;
	wire [0:0] ejection_channels_403__bench;
	wire [0:0] ejection_channels_402__bench;
	wire [0:0] ejection_channels_401__bench;
	wire [0:0] ejection_channels_400__bench;
	wire [0:0] ejection_channels_399__bench;
	wire [0:0] ejection_channels_398__bench;
	wire [0:0] ejection_channels_397__bench;
	wire [0:0] ejection_channels_396__bench;
	wire [0:0] ejection_channels_395__bench;
	wire [0:0] ejection_channels_394__bench;
	wire [0:0] ejection_channels_393__bench;
	wire [0:0] ejection_channels_392__bench;
	wire [0:0] ejection_channels_391__bench;
	wire [0:0] ejection_channels_390__bench;
	wire [0:0] ejection_channels_389__bench;
	wire [0:0] ejection_channels_388__bench;
	wire [0:0] ejection_channels_387__bench;
	wire [0:0] ejection_channels_386__bench;
	wire [0:0] ejection_channels_385__bench;
	wire [0:0] ejection_channels_384__bench;
	wire [0:0] ejection_channels_383__bench;
	wire [0:0] ejection_channels_382__bench;
	wire [0:0] ejection_channels_381__bench;
	wire [0:0] ejection_channels_380__bench;
	wire [0:0] ejection_channels_379__bench;
	wire [0:0] ejection_channels_378__bench;
	wire [0:0] ejection_channels_377__bench;
	wire [0:0] ejection_channels_376__bench;
	wire [0:0] ejection_channels_375__bench;
	wire [0:0] ejection_channels_374__bench;
	wire [0:0] ejection_channels_373__bench;
	wire [0:0] ejection_channels_372__bench;
	wire [0:0] ejection_channels_371__bench;
	wire [0:0] ejection_channels_370__bench;
	wire [0:0] ejection_channels_369__bench;
	wire [0:0] ejection_channels_368__bench;
	wire [0:0] ejection_channels_367__bench;
	wire [0:0] ejection_channels_366__bench;
	wire [0:0] ejection_channels_365__bench;
	wire [0:0] ejection_channels_364__bench;
	wire [0:0] ejection_channels_363__bench;
	wire [0:0] ejection_channels_362__bench;
	wire [0:0] ejection_channels_361__bench;
	wire [0:0] ejection_channels_360__bench;
	wire [0:0] ejection_channels_359__bench;
	wire [0:0] ejection_channels_358__bench;
	wire [0:0] ejection_channels_357__bench;
	wire [0:0] ejection_channels_356__bench;
	wire [0:0] ejection_channels_355__bench;
	wire [0:0] ejection_channels_354__bench;
	wire [0:0] ejection_channels_353__bench;
	wire [0:0] ejection_channels_352__bench;
	wire [0:0] ejection_channels_351__bench;
	wire [0:0] ejection_channels_350__bench;
	wire [0:0] ejection_channels_349__bench;
	wire [0:0] ejection_channels_348__bench;
	wire [0:0] ejection_channels_347__bench;
	wire [0:0] ejection_channels_346__bench;
	wire [0:0] ejection_channels_345__bench;
	wire [0:0] ejection_channels_344__bench;
	wire [0:0] ejection_channels_343__bench;
	wire [0:0] ejection_channels_342__bench;
	wire [0:0] ejection_channels_341__bench;
	wire [0:0] ejection_channels_340__bench;
	wire [0:0] ejection_channels_339__bench;
	wire [0:0] ejection_channels_338__bench;
	wire [0:0] ejection_channels_337__bench;
	wire [0:0] ejection_channels_336__bench;
	wire [0:0] ejection_channels_335__bench;
	wire [0:0] ejection_channels_334__bench;
	wire [0:0] ejection_channels_333__bench;
	wire [0:0] ejection_channels_332__bench;
	wire [0:0] ejection_channels_331__bench;
	wire [0:0] ejection_channels_330__bench;
	wire [0:0] ejection_channels_329__bench;
	wire [0:0] ejection_channels_328__bench;
	wire [0:0] ejection_channels_327__bench;
	wire [0:0] ejection_channels_326__bench;
	wire [0:0] ejection_channels_325__bench;
	wire [0:0] ejection_channels_324__bench;
	wire [0:0] ejection_channels_323__bench;
	wire [0:0] ejection_channels_322__bench;
	wire [0:0] ejection_channels_321__bench;
	wire [0:0] ejection_channels_320__bench;
	wire [0:0] ejection_channels_319__bench;
	wire [0:0] ejection_channels_318__bench;
	wire [0:0] ejection_channels_317__bench;
	wire [0:0] ejection_channels_316__bench;
	wire [0:0] ejection_channels_315__bench;
	wire [0:0] ejection_channels_314__bench;
	wire [0:0] ejection_channels_313__bench;
	wire [0:0] ejection_channels_312__bench;
	wire [0:0] ejection_channels_311__bench;
	wire [0:0] ejection_channels_310__bench;
	wire [0:0] ejection_channels_309__bench;
	wire [0:0] ejection_channels_308__bench;
	wire [0:0] ejection_channels_307__bench;
	wire [0:0] ejection_channels_306__bench;
	wire [0:0] ejection_channels_305__bench;
	wire [0:0] ejection_channels_304__bench;
	wire [0:0] ejection_channels_303__bench;
	wire [0:0] ejection_channels_302__bench;
	wire [0:0] ejection_channels_301__bench;
	wire [0:0] ejection_channels_300__bench;
	wire [0:0] ejection_channels_299__bench;
	wire [0:0] ejection_channels_298__bench;
	wire [0:0] ejection_channels_297__bench;
	wire [0:0] ejection_channels_296__bench;
	wire [0:0] ejection_channels_295__bench;
	wire [0:0] ejection_channels_294__bench;
	wire [0:0] ejection_channels_293__bench;
	wire [0:0] ejection_channels_292__bench;
	wire [0:0] ejection_channels_291__bench;
	wire [0:0] ejection_channels_290__bench;
	wire [0:0] ejection_channels_289__bench;
	wire [0:0] ejection_channels_288__bench;
	wire [0:0] ejection_channels_287__bench;
	wire [0:0] ejection_channels_286__bench;
	wire [0:0] ejection_channels_285__bench;
	wire [0:0] ejection_channels_284__bench;
	wire [0:0] ejection_channels_283__bench;
	wire [0:0] ejection_channels_282__bench;
	wire [0:0] ejection_channels_281__bench;
	wire [0:0] ejection_channels_280__bench;
	wire [0:0] ejection_channels_279__bench;
	wire [0:0] ejection_channels_278__bench;
	wire [0:0] ejection_channels_277__bench;
	wire [0:0] ejection_channels_276__bench;
	wire [0:0] ejection_channels_275__bench;
	wire [0:0] ejection_channels_274__bench;
	wire [0:0] ejection_channels_273__bench;
	wire [0:0] ejection_channels_272__bench;
	wire [0:0] ejection_channels_271__bench;
	wire [0:0] ejection_channels_270__bench;
	wire [0:0] ejection_channels_269__bench;
	wire [0:0] ejection_channels_268__bench;
	wire [0:0] ejection_channels_267__bench;
	wire [0:0] ejection_channels_266__bench;
	wire [0:0] ejection_channels_265__bench;
	wire [0:0] ejection_channels_264__bench;
	wire [0:0] ejection_channels_263__bench;
	wire [0:0] ejection_channels_262__bench;
	wire [0:0] ejection_channels_261__bench;
	wire [0:0] ejection_channels_260__bench;
	wire [0:0] ejection_channels_259__bench;
	wire [0:0] ejection_channels_258__bench;
	wire [0:0] ejection_channels_257__bench;
	wire [0:0] ejection_channels_256__bench;
	wire [0:0] ejection_channels_255__bench;
	wire [0:0] ejection_channels_254__bench;
	wire [0:0] ejection_channels_253__bench;
	wire [0:0] ejection_channels_252__bench;
	wire [0:0] ejection_channels_251__bench;
	wire [0:0] ejection_channels_250__bench;
	wire [0:0] ejection_channels_249__bench;
	wire [0:0] ejection_channels_248__bench;
	wire [0:0] ejection_channels_247__bench;
	wire [0:0] ejection_channels_246__bench;
	wire [0:0] ejection_channels_245__bench;
	wire [0:0] ejection_channels_244__bench;
	wire [0:0] ejection_channels_243__bench;
	wire [0:0] ejection_channels_242__bench;
	wire [0:0] ejection_channels_241__bench;
	wire [0:0] ejection_channels_240__bench;
	wire [0:0] ejection_channels_239__bench;
	wire [0:0] ejection_channels_238__bench;
	wire [0:0] ejection_channels_237__bench;
	wire [0:0] ejection_channels_236__bench;
	wire [0:0] ejection_channels_235__bench;
	wire [0:0] ejection_channels_234__bench;
	wire [0:0] ejection_channels_233__bench;
	wire [0:0] ejection_channels_232__bench;
	wire [0:0] ejection_channels_231__bench;
	wire [0:0] ejection_channels_230__bench;
	wire [0:0] ejection_channels_229__bench;
	wire [0:0] ejection_channels_228__bench;
	wire [0:0] ejection_channels_227__bench;
	wire [0:0] ejection_channels_226__bench;
	wire [0:0] ejection_channels_225__bench;
	wire [0:0] ejection_channels_224__bench;
	wire [0:0] ejection_channels_223__bench;
	wire [0:0] ejection_channels_222__bench;
	wire [0:0] ejection_channels_221__bench;
	wire [0:0] ejection_channels_220__bench;
	wire [0:0] ejection_channels_219__bench;
	wire [0:0] ejection_channels_218__bench;
	wire [0:0] ejection_channels_217__bench;
	wire [0:0] ejection_channels_216__bench;
	wire [0:0] ejection_channels_215__bench;
	wire [0:0] ejection_channels_214__bench;
	wire [0:0] ejection_channels_213__bench;
	wire [0:0] ejection_channels_212__bench;
	wire [0:0] ejection_channels_211__bench;
	wire [0:0] ejection_channels_210__bench;
	wire [0:0] ejection_channels_209__bench;
	wire [0:0] ejection_channels_208__bench;
	wire [0:0] ejection_channels_207__bench;
	wire [0:0] ejection_channels_206__bench;
	wire [0:0] ejection_channels_205__bench;
	wire [0:0] ejection_channels_204__bench;
	wire [0:0] ejection_channels_203__bench;
	wire [0:0] ejection_channels_202__bench;
	wire [0:0] ejection_channels_201__bench;
	wire [0:0] ejection_channels_200__bench;
	wire [0:0] ejection_channels_199__bench;
	wire [0:0] ejection_channels_198__bench;
	wire [0:0] ejection_channels_197__bench;
	wire [0:0] ejection_channels_196__bench;
	wire [0:0] ejection_channels_195__bench;
	wire [0:0] ejection_channels_194__bench;
	wire [0:0] ejection_channels_193__bench;
	wire [0:0] ejection_channels_192__bench;
	wire [0:0] ejection_channels_191__bench;
	wire [0:0] ejection_channels_190__bench;
	wire [0:0] ejection_channels_189__bench;
	wire [0:0] ejection_channels_188__bench;
	wire [0:0] ejection_channels_187__bench;
	wire [0:0] ejection_channels_186__bench;
	wire [0:0] ejection_channels_185__bench;
	wire [0:0] ejection_channels_184__bench;
	wire [0:0] ejection_channels_183__bench;
	wire [0:0] ejection_channels_182__bench;
	wire [0:0] ejection_channels_181__bench;
	wire [0:0] ejection_channels_180__bench;
	wire [0:0] ejection_channels_179__bench;
	wire [0:0] ejection_channels_178__bench;
	wire [0:0] ejection_channels_177__bench;
	wire [0:0] ejection_channels_176__bench;
	wire [0:0] ejection_channels_175__bench;
	wire [0:0] ejection_channels_174__bench;
	wire [0:0] ejection_channels_173__bench;
	wire [0:0] ejection_channels_172__bench;
	wire [0:0] ejection_channels_171__bench;
	wire [0:0] ejection_channels_170__bench;
	wire [0:0] ejection_channels_169__bench;
	wire [0:0] ejection_channels_168__bench;
	wire [0:0] ejection_channels_167__bench;
	wire [0:0] ejection_channels_166__bench;
	wire [0:0] ejection_channels_165__bench;
	wire [0:0] ejection_channels_164__bench;
	wire [0:0] ejection_channels_163__bench;
	wire [0:0] ejection_channels_162__bench;
	wire [0:0] ejection_channels_161__bench;
	wire [0:0] ejection_channels_160__bench;
	wire [0:0] ejection_channels_159__bench;
	wire [0:0] ejection_channels_158__bench;
	wire [0:0] ejection_channels_157__bench;
	wire [0:0] ejection_channels_156__bench;
	wire [0:0] ejection_channels_155__bench;
	wire [0:0] ejection_channels_154__bench;
	wire [0:0] ejection_channels_153__bench;
	wire [0:0] ejection_channels_152__bench;
	wire [0:0] ejection_channels_151__bench;
	wire [0:0] ejection_channels_150__bench;
	wire [0:0] ejection_channels_149__bench;
	wire [0:0] ejection_channels_148__bench;
	wire [0:0] ejection_channels_147__bench;
	wire [0:0] ejection_channels_146__bench;
	wire [0:0] ejection_channels_145__bench;
	wire [0:0] ejection_channels_144__bench;
	wire [0:0] ejection_channels_143__bench;
	wire [0:0] ejection_channels_142__bench;
	wire [0:0] ejection_channels_141__bench;
	wire [0:0] ejection_channels_140__bench;
	wire [0:0] ejection_channels_139__bench;
	wire [0:0] ejection_channels_138__bench;
	wire [0:0] ejection_channels_137__bench;
	wire [0:0] ejection_channels_136__bench;
	wire [0:0] ejection_channels_135__bench;
	wire [0:0] ejection_channels_134__bench;
	wire [0:0] ejection_channels_133__bench;
	wire [0:0] ejection_channels_132__bench;
	wire [0:0] ejection_channels_131__bench;
	wire [0:0] ejection_channels_130__bench;
	wire [0:0] ejection_channels_129__bench;
	wire [0:0] ejection_channels_128__bench;
	wire [0:0] ejection_channels_127__bench;
	wire [0:0] ejection_channels_126__bench;
	wire [0:0] ejection_channels_125__bench;
	wire [0:0] ejection_channels_124__bench;
	wire [0:0] ejection_channels_123__bench;
	wire [0:0] ejection_channels_122__bench;
	wire [0:0] ejection_channels_121__bench;
	wire [0:0] ejection_channels_120__bench;
	wire [0:0] ejection_channels_119__bench;
	wire [0:0] ejection_channels_118__bench;
	wire [0:0] ejection_channels_117__bench;
	wire [0:0] ejection_channels_116__bench;
	wire [0:0] ejection_channels_115__bench;
	wire [0:0] ejection_channels_114__bench;
	wire [0:0] ejection_channels_113__bench;
	wire [0:0] ejection_channels_112__bench;
	wire [0:0] ejection_channels_111__bench;
	wire [0:0] ejection_channels_110__bench;
	wire [0:0] ejection_channels_109__bench;
	wire [0:0] ejection_channels_108__bench;
	wire [0:0] ejection_channels_107__bench;
	wire [0:0] ejection_channels_106__bench;
	wire [0:0] ejection_channels_105__bench;
	wire [0:0] ejection_channels_104__bench;
	wire [0:0] ejection_channels_103__bench;
	wire [0:0] ejection_channels_102__bench;
	wire [0:0] ejection_channels_101__bench;
	wire [0:0] ejection_channels_100__bench;
	wire [0:0] ejection_channels_99__bench;
	wire [0:0] ejection_channels_98__bench;
	wire [0:0] ejection_channels_97__bench;
	wire [0:0] ejection_channels_96__bench;
	wire [0:0] ejection_channels_95__bench;
	wire [0:0] ejection_channels_94__bench;
	wire [0:0] ejection_channels_93__bench;
	wire [0:0] ejection_channels_92__bench;
	wire [0:0] ejection_channels_91__bench;
	wire [0:0] ejection_channels_90__bench;
	wire [0:0] ejection_channels_89__bench;
	wire [0:0] ejection_channels_88__bench;
	wire [0:0] ejection_channels_87__bench;
	wire [0:0] ejection_channels_86__bench;
	wire [0:0] ejection_channels_85__bench;
	wire [0:0] ejection_channels_84__bench;
	wire [0:0] ejection_channels_83__bench;
	wire [0:0] ejection_channels_82__bench;
	wire [0:0] ejection_channels_81__bench;
	wire [0:0] ejection_channels_80__bench;
	wire [0:0] ejection_channels_79__bench;
	wire [0:0] ejection_channels_78__bench;
	wire [0:0] ejection_channels_77__bench;
	wire [0:0] ejection_channels_76__bench;
	wire [0:0] ejection_channels_75__bench;
	wire [0:0] ejection_channels_74__bench;
	wire [0:0] ejection_channels_73__bench;
	wire [0:0] ejection_channels_72__bench;
	wire [0:0] ejection_channels_71__bench;
	wire [0:0] ejection_channels_70__bench;
	wire [0:0] ejection_channels_69__bench;
	wire [0:0] ejection_channels_68__bench;
	wire [0:0] ejection_channels_67__bench;
	wire [0:0] ejection_channels_66__bench;
	wire [0:0] ejection_channels_65__bench;
	wire [0:0] ejection_channels_64__bench;
	wire [0:0] ejection_channels_63__bench;
	wire [0:0] ejection_channels_62__bench;
	wire [0:0] ejection_channels_61__bench;
	wire [0:0] ejection_channels_60__bench;
	wire [0:0] ejection_channels_59__bench;
	wire [0:0] ejection_channels_58__bench;
	wire [0:0] ejection_channels_57__bench;
	wire [0:0] ejection_channels_56__bench;
	wire [0:0] ejection_channels_55__bench;
	wire [0:0] ejection_channels_54__bench;
	wire [0:0] ejection_channels_53__bench;
	wire [0:0] ejection_channels_52__bench;
	wire [0:0] ejection_channels_51__bench;
	wire [0:0] ejection_channels_50__bench;
	wire [0:0] ejection_channels_49__bench;
	wire [0:0] ejection_channels_48__bench;
	wire [0:0] ejection_channels_47__bench;
	wire [0:0] ejection_channels_46__bench;
	wire [0:0] ejection_channels_45__bench;
	wire [0:0] ejection_channels_44__bench;
	wire [0:0] ejection_channels_43__bench;
	wire [0:0] ejection_channels_42__bench;
	wire [0:0] ejection_channels_41__bench;
	wire [0:0] ejection_channels_40__bench;
	wire [0:0] ejection_channels_39__bench;
	wire [0:0] ejection_channels_38__bench;
	wire [0:0] ejection_channels_37__bench;
	wire [0:0] ejection_channels_36__bench;
	wire [0:0] ejection_channels_35__bench;
	wire [0:0] ejection_channels_34__bench;
	wire [0:0] ejection_channels_33__bench;
	wire [0:0] ejection_channels_32__bench;
	wire [0:0] ejection_channels_31__bench;
	wire [0:0] ejection_channels_30__bench;
	wire [0:0] ejection_channels_29__bench;
	wire [0:0] ejection_channels_28__bench;
	wire [0:0] ejection_channels_27__bench;
	wire [0:0] ejection_channels_26__bench;
	wire [0:0] ejection_channels_25__bench;
	wire [0:0] ejection_channels_24__bench;
	wire [0:0] ejection_channels_23__bench;
	wire [0:0] ejection_channels_22__bench;
	wire [0:0] ejection_channels_21__bench;
	wire [0:0] ejection_channels_20__bench;
	wire [0:0] ejection_channels_19__bench;
	wire [0:0] ejection_channels_18__bench;
	wire [0:0] ejection_channels_17__bench;
	wire [0:0] ejection_channels_16__bench;
	wire [0:0] ejection_channels_15__bench;
	wire [0:0] ejection_channels_14__bench;
	wire [0:0] ejection_channels_13__bench;
	wire [0:0] ejection_channels_12__bench;
	wire [0:0] ejection_channels_11__bench;
	wire [0:0] ejection_channels_10__bench;
	wire [0:0] ejection_channels_9__bench;
	wire [0:0] ejection_channels_8__bench;
	wire [0:0] ejection_channels_7__bench;
	wire [0:0] ejection_channels_6__bench;
	wire [0:0] ejection_channels_5__bench;
	wire [0:0] ejection_channels_4__bench;
	wire [0:0] ejection_channels_3__bench;
	wire [0:0] ejection_channels_2__bench;
	wire [0:0] ejection_channels_1__bench;
	wire [0:0] ejection_channels_0__bench;
	wire [0:0] rtr_error_8__bench;
	wire [0:0] rtr_error_7__bench;
	wire [0:0] rtr_error_6__bench;
	wire [0:0] rtr_error_5__bench;
	wire [0:0] rtr_error_4__bench;
	wire [0:0] rtr_error_3__bench;
	wire [0:0] rtr_error_2__bench;
	wire [0:0] rtr_error_1__bench;
	wire [0:0] rtr_error_0__bench;

// ----- Output vectors checking flags -------
	reg [0:0] injection_flow_ctrl_26__flag;
	reg [0:0] injection_flow_ctrl_25__flag;
	reg [0:0] injection_flow_ctrl_24__flag;
	reg [0:0] injection_flow_ctrl_23__flag;
	reg [0:0] injection_flow_ctrl_22__flag;
	reg [0:0] injection_flow_ctrl_21__flag;
	reg [0:0] injection_flow_ctrl_20__flag;
	reg [0:0] injection_flow_ctrl_19__flag;
	reg [0:0] injection_flow_ctrl_18__flag;
	reg [0:0] injection_flow_ctrl_17__flag;
	reg [0:0] injection_flow_ctrl_16__flag;
	reg [0:0] injection_flow_ctrl_15__flag;
	reg [0:0] injection_flow_ctrl_14__flag;
	reg [0:0] injection_flow_ctrl_13__flag;
	reg [0:0] injection_flow_ctrl_12__flag;
	reg [0:0] injection_flow_ctrl_11__flag;
	reg [0:0] injection_flow_ctrl_10__flag;
	reg [0:0] injection_flow_ctrl_9__flag;
	reg [0:0] injection_flow_ctrl_8__flag;
	reg [0:0] injection_flow_ctrl_7__flag;
	reg [0:0] injection_flow_ctrl_6__flag;
	reg [0:0] injection_flow_ctrl_5__flag;
	reg [0:0] injection_flow_ctrl_4__flag;
	reg [0:0] injection_flow_ctrl_3__flag;
	reg [0:0] injection_flow_ctrl_2__flag;
	reg [0:0] injection_flow_ctrl_1__flag;
	reg [0:0] injection_flow_ctrl_0__flag;
	reg [0:0] ejection_channels_629__flag;
	reg [0:0] ejection_channels_628__flag;
	reg [0:0] ejection_channels_627__flag;
	reg [0:0] ejection_channels_626__flag;
	reg [0:0] ejection_channels_625__flag;
	reg [0:0] ejection_channels_624__flag;
	reg [0:0] ejection_channels_623__flag;
	reg [0:0] ejection_channels_622__flag;
	reg [0:0] ejection_channels_621__flag;
	reg [0:0] ejection_channels_620__flag;
	reg [0:0] ejection_channels_619__flag;
	reg [0:0] ejection_channels_618__flag;
	reg [0:0] ejection_channels_617__flag;
	reg [0:0] ejection_channels_616__flag;
	reg [0:0] ejection_channels_615__flag;
	reg [0:0] ejection_channels_614__flag;
	reg [0:0] ejection_channels_613__flag;
	reg [0:0] ejection_channels_612__flag;
	reg [0:0] ejection_channels_611__flag;
	reg [0:0] ejection_channels_610__flag;
	reg [0:0] ejection_channels_609__flag;
	reg [0:0] ejection_channels_608__flag;
	reg [0:0] ejection_channels_607__flag;
	reg [0:0] ejection_channels_606__flag;
	reg [0:0] ejection_channels_605__flag;
	reg [0:0] ejection_channels_604__flag;
	reg [0:0] ejection_channels_603__flag;
	reg [0:0] ejection_channels_602__flag;
	reg [0:0] ejection_channels_601__flag;
	reg [0:0] ejection_channels_600__flag;
	reg [0:0] ejection_channels_599__flag;
	reg [0:0] ejection_channels_598__flag;
	reg [0:0] ejection_channels_597__flag;
	reg [0:0] ejection_channels_596__flag;
	reg [0:0] ejection_channels_595__flag;
	reg [0:0] ejection_channels_594__flag;
	reg [0:0] ejection_channels_593__flag;
	reg [0:0] ejection_channels_592__flag;
	reg [0:0] ejection_channels_591__flag;
	reg [0:0] ejection_channels_590__flag;
	reg [0:0] ejection_channels_589__flag;
	reg [0:0] ejection_channels_588__flag;
	reg [0:0] ejection_channels_587__flag;
	reg [0:0] ejection_channels_586__flag;
	reg [0:0] ejection_channels_585__flag;
	reg [0:0] ejection_channels_584__flag;
	reg [0:0] ejection_channels_583__flag;
	reg [0:0] ejection_channels_582__flag;
	reg [0:0] ejection_channels_581__flag;
	reg [0:0] ejection_channels_580__flag;
	reg [0:0] ejection_channels_579__flag;
	reg [0:0] ejection_channels_578__flag;
	reg [0:0] ejection_channels_577__flag;
	reg [0:0] ejection_channels_576__flag;
	reg [0:0] ejection_channels_575__flag;
	reg [0:0] ejection_channels_574__flag;
	reg [0:0] ejection_channels_573__flag;
	reg [0:0] ejection_channels_572__flag;
	reg [0:0] ejection_channels_571__flag;
	reg [0:0] ejection_channels_570__flag;
	reg [0:0] ejection_channels_569__flag;
	reg [0:0] ejection_channels_568__flag;
	reg [0:0] ejection_channels_567__flag;
	reg [0:0] ejection_channels_566__flag;
	reg [0:0] ejection_channels_565__flag;
	reg [0:0] ejection_channels_564__flag;
	reg [0:0] ejection_channels_563__flag;
	reg [0:0] ejection_channels_562__flag;
	reg [0:0] ejection_channels_561__flag;
	reg [0:0] ejection_channels_560__flag;
	reg [0:0] ejection_channels_559__flag;
	reg [0:0] ejection_channels_558__flag;
	reg [0:0] ejection_channels_557__flag;
	reg [0:0] ejection_channels_556__flag;
	reg [0:0] ejection_channels_555__flag;
	reg [0:0] ejection_channels_554__flag;
	reg [0:0] ejection_channels_553__flag;
	reg [0:0] ejection_channels_552__flag;
	reg [0:0] ejection_channels_551__flag;
	reg [0:0] ejection_channels_550__flag;
	reg [0:0] ejection_channels_549__flag;
	reg [0:0] ejection_channels_548__flag;
	reg [0:0] ejection_channels_547__flag;
	reg [0:0] ejection_channels_546__flag;
	reg [0:0] ejection_channels_545__flag;
	reg [0:0] ejection_channels_544__flag;
	reg [0:0] ejection_channels_543__flag;
	reg [0:0] ejection_channels_542__flag;
	reg [0:0] ejection_channels_541__flag;
	reg [0:0] ejection_channels_540__flag;
	reg [0:0] ejection_channels_539__flag;
	reg [0:0] ejection_channels_538__flag;
	reg [0:0] ejection_channels_537__flag;
	reg [0:0] ejection_channels_536__flag;
	reg [0:0] ejection_channels_535__flag;
	reg [0:0] ejection_channels_534__flag;
	reg [0:0] ejection_channels_533__flag;
	reg [0:0] ejection_channels_532__flag;
	reg [0:0] ejection_channels_531__flag;
	reg [0:0] ejection_channels_530__flag;
	reg [0:0] ejection_channels_529__flag;
	reg [0:0] ejection_channels_528__flag;
	reg [0:0] ejection_channels_527__flag;
	reg [0:0] ejection_channels_526__flag;
	reg [0:0] ejection_channels_525__flag;
	reg [0:0] ejection_channels_524__flag;
	reg [0:0] ejection_channels_523__flag;
	reg [0:0] ejection_channels_522__flag;
	reg [0:0] ejection_channels_521__flag;
	reg [0:0] ejection_channels_520__flag;
	reg [0:0] ejection_channels_519__flag;
	reg [0:0] ejection_channels_518__flag;
	reg [0:0] ejection_channels_517__flag;
	reg [0:0] ejection_channels_516__flag;
	reg [0:0] ejection_channels_515__flag;
	reg [0:0] ejection_channels_514__flag;
	reg [0:0] ejection_channels_513__flag;
	reg [0:0] ejection_channels_512__flag;
	reg [0:0] ejection_channels_511__flag;
	reg [0:0] ejection_channels_510__flag;
	reg [0:0] ejection_channels_509__flag;
	reg [0:0] ejection_channels_508__flag;
	reg [0:0] ejection_channels_507__flag;
	reg [0:0] ejection_channels_506__flag;
	reg [0:0] ejection_channels_505__flag;
	reg [0:0] ejection_channels_504__flag;
	reg [0:0] ejection_channels_503__flag;
	reg [0:0] ejection_channels_502__flag;
	reg [0:0] ejection_channels_501__flag;
	reg [0:0] ejection_channels_500__flag;
	reg [0:0] ejection_channels_499__flag;
	reg [0:0] ejection_channels_498__flag;
	reg [0:0] ejection_channels_497__flag;
	reg [0:0] ejection_channels_496__flag;
	reg [0:0] ejection_channels_495__flag;
	reg [0:0] ejection_channels_494__flag;
	reg [0:0] ejection_channels_493__flag;
	reg [0:0] ejection_channels_492__flag;
	reg [0:0] ejection_channels_491__flag;
	reg [0:0] ejection_channels_490__flag;
	reg [0:0] ejection_channels_489__flag;
	reg [0:0] ejection_channels_488__flag;
	reg [0:0] ejection_channels_487__flag;
	reg [0:0] ejection_channels_486__flag;
	reg [0:0] ejection_channels_485__flag;
	reg [0:0] ejection_channels_484__flag;
	reg [0:0] ejection_channels_483__flag;
	reg [0:0] ejection_channels_482__flag;
	reg [0:0] ejection_channels_481__flag;
	reg [0:0] ejection_channels_480__flag;
	reg [0:0] ejection_channels_479__flag;
	reg [0:0] ejection_channels_478__flag;
	reg [0:0] ejection_channels_477__flag;
	reg [0:0] ejection_channels_476__flag;
	reg [0:0] ejection_channels_475__flag;
	reg [0:0] ejection_channels_474__flag;
	reg [0:0] ejection_channels_473__flag;
	reg [0:0] ejection_channels_472__flag;
	reg [0:0] ejection_channels_471__flag;
	reg [0:0] ejection_channels_470__flag;
	reg [0:0] ejection_channels_469__flag;
	reg [0:0] ejection_channels_468__flag;
	reg [0:0] ejection_channels_467__flag;
	reg [0:0] ejection_channels_466__flag;
	reg [0:0] ejection_channels_465__flag;
	reg [0:0] ejection_channels_464__flag;
	reg [0:0] ejection_channels_463__flag;
	reg [0:0] ejection_channels_462__flag;
	reg [0:0] ejection_channels_461__flag;
	reg [0:0] ejection_channels_460__flag;
	reg [0:0] ejection_channels_459__flag;
	reg [0:0] ejection_channels_458__flag;
	reg [0:0] ejection_channels_457__flag;
	reg [0:0] ejection_channels_456__flag;
	reg [0:0] ejection_channels_455__flag;
	reg [0:0] ejection_channels_454__flag;
	reg [0:0] ejection_channels_453__flag;
	reg [0:0] ejection_channels_452__flag;
	reg [0:0] ejection_channels_451__flag;
	reg [0:0] ejection_channels_450__flag;
	reg [0:0] ejection_channels_449__flag;
	reg [0:0] ejection_channels_448__flag;
	reg [0:0] ejection_channels_447__flag;
	reg [0:0] ejection_channels_446__flag;
	reg [0:0] ejection_channels_445__flag;
	reg [0:0] ejection_channels_444__flag;
	reg [0:0] ejection_channels_443__flag;
	reg [0:0] ejection_channels_442__flag;
	reg [0:0] ejection_channels_441__flag;
	reg [0:0] ejection_channels_440__flag;
	reg [0:0] ejection_channels_439__flag;
	reg [0:0] ejection_channels_438__flag;
	reg [0:0] ejection_channels_437__flag;
	reg [0:0] ejection_channels_436__flag;
	reg [0:0] ejection_channels_435__flag;
	reg [0:0] ejection_channels_434__flag;
	reg [0:0] ejection_channels_433__flag;
	reg [0:0] ejection_channels_432__flag;
	reg [0:0] ejection_channels_431__flag;
	reg [0:0] ejection_channels_430__flag;
	reg [0:0] ejection_channels_429__flag;
	reg [0:0] ejection_channels_428__flag;
	reg [0:0] ejection_channels_427__flag;
	reg [0:0] ejection_channels_426__flag;
	reg [0:0] ejection_channels_425__flag;
	reg [0:0] ejection_channels_424__flag;
	reg [0:0] ejection_channels_423__flag;
	reg [0:0] ejection_channels_422__flag;
	reg [0:0] ejection_channels_421__flag;
	reg [0:0] ejection_channels_420__flag;
	reg [0:0] ejection_channels_419__flag;
	reg [0:0] ejection_channels_418__flag;
	reg [0:0] ejection_channels_417__flag;
	reg [0:0] ejection_channels_416__flag;
	reg [0:0] ejection_channels_415__flag;
	reg [0:0] ejection_channels_414__flag;
	reg [0:0] ejection_channels_413__flag;
	reg [0:0] ejection_channels_412__flag;
	reg [0:0] ejection_channels_411__flag;
	reg [0:0] ejection_channels_410__flag;
	reg [0:0] ejection_channels_409__flag;
	reg [0:0] ejection_channels_408__flag;
	reg [0:0] ejection_channels_407__flag;
	reg [0:0] ejection_channels_406__flag;
	reg [0:0] ejection_channels_405__flag;
	reg [0:0] ejection_channels_404__flag;
	reg [0:0] ejection_channels_403__flag;
	reg [0:0] ejection_channels_402__flag;
	reg [0:0] ejection_channels_401__flag;
	reg [0:0] ejection_channels_400__flag;
	reg [0:0] ejection_channels_399__flag;
	reg [0:0] ejection_channels_398__flag;
	reg [0:0] ejection_channels_397__flag;
	reg [0:0] ejection_channels_396__flag;
	reg [0:0] ejection_channels_395__flag;
	reg [0:0] ejection_channels_394__flag;
	reg [0:0] ejection_channels_393__flag;
	reg [0:0] ejection_channels_392__flag;
	reg [0:0] ejection_channels_391__flag;
	reg [0:0] ejection_channels_390__flag;
	reg [0:0] ejection_channels_389__flag;
	reg [0:0] ejection_channels_388__flag;
	reg [0:0] ejection_channels_387__flag;
	reg [0:0] ejection_channels_386__flag;
	reg [0:0] ejection_channels_385__flag;
	reg [0:0] ejection_channels_384__flag;
	reg [0:0] ejection_channels_383__flag;
	reg [0:0] ejection_channels_382__flag;
	reg [0:0] ejection_channels_381__flag;
	reg [0:0] ejection_channels_380__flag;
	reg [0:0] ejection_channels_379__flag;
	reg [0:0] ejection_channels_378__flag;
	reg [0:0] ejection_channels_377__flag;
	reg [0:0] ejection_channels_376__flag;
	reg [0:0] ejection_channels_375__flag;
	reg [0:0] ejection_channels_374__flag;
	reg [0:0] ejection_channels_373__flag;
	reg [0:0] ejection_channels_372__flag;
	reg [0:0] ejection_channels_371__flag;
	reg [0:0] ejection_channels_370__flag;
	reg [0:0] ejection_channels_369__flag;
	reg [0:0] ejection_channels_368__flag;
	reg [0:0] ejection_channels_367__flag;
	reg [0:0] ejection_channels_366__flag;
	reg [0:0] ejection_channels_365__flag;
	reg [0:0] ejection_channels_364__flag;
	reg [0:0] ejection_channels_363__flag;
	reg [0:0] ejection_channels_362__flag;
	reg [0:0] ejection_channels_361__flag;
	reg [0:0] ejection_channels_360__flag;
	reg [0:0] ejection_channels_359__flag;
	reg [0:0] ejection_channels_358__flag;
	reg [0:0] ejection_channels_357__flag;
	reg [0:0] ejection_channels_356__flag;
	reg [0:0] ejection_channels_355__flag;
	reg [0:0] ejection_channels_354__flag;
	reg [0:0] ejection_channels_353__flag;
	reg [0:0] ejection_channels_352__flag;
	reg [0:0] ejection_channels_351__flag;
	reg [0:0] ejection_channels_350__flag;
	reg [0:0] ejection_channels_349__flag;
	reg [0:0] ejection_channels_348__flag;
	reg [0:0] ejection_channels_347__flag;
	reg [0:0] ejection_channels_346__flag;
	reg [0:0] ejection_channels_345__flag;
	reg [0:0] ejection_channels_344__flag;
	reg [0:0] ejection_channels_343__flag;
	reg [0:0] ejection_channels_342__flag;
	reg [0:0] ejection_channels_341__flag;
	reg [0:0] ejection_channels_340__flag;
	reg [0:0] ejection_channels_339__flag;
	reg [0:0] ejection_channels_338__flag;
	reg [0:0] ejection_channels_337__flag;
	reg [0:0] ejection_channels_336__flag;
	reg [0:0] ejection_channels_335__flag;
	reg [0:0] ejection_channels_334__flag;
	reg [0:0] ejection_channels_333__flag;
	reg [0:0] ejection_channels_332__flag;
	reg [0:0] ejection_channels_331__flag;
	reg [0:0] ejection_channels_330__flag;
	reg [0:0] ejection_channels_329__flag;
	reg [0:0] ejection_channels_328__flag;
	reg [0:0] ejection_channels_327__flag;
	reg [0:0] ejection_channels_326__flag;
	reg [0:0] ejection_channels_325__flag;
	reg [0:0] ejection_channels_324__flag;
	reg [0:0] ejection_channels_323__flag;
	reg [0:0] ejection_channels_322__flag;
	reg [0:0] ejection_channels_321__flag;
	reg [0:0] ejection_channels_320__flag;
	reg [0:0] ejection_channels_319__flag;
	reg [0:0] ejection_channels_318__flag;
	reg [0:0] ejection_channels_317__flag;
	reg [0:0] ejection_channels_316__flag;
	reg [0:0] ejection_channels_315__flag;
	reg [0:0] ejection_channels_314__flag;
	reg [0:0] ejection_channels_313__flag;
	reg [0:0] ejection_channels_312__flag;
	reg [0:0] ejection_channels_311__flag;
	reg [0:0] ejection_channels_310__flag;
	reg [0:0] ejection_channels_309__flag;
	reg [0:0] ejection_channels_308__flag;
	reg [0:0] ejection_channels_307__flag;
	reg [0:0] ejection_channels_306__flag;
	reg [0:0] ejection_channels_305__flag;
	reg [0:0] ejection_channels_304__flag;
	reg [0:0] ejection_channels_303__flag;
	reg [0:0] ejection_channels_302__flag;
	reg [0:0] ejection_channels_301__flag;
	reg [0:0] ejection_channels_300__flag;
	reg [0:0] ejection_channels_299__flag;
	reg [0:0] ejection_channels_298__flag;
	reg [0:0] ejection_channels_297__flag;
	reg [0:0] ejection_channels_296__flag;
	reg [0:0] ejection_channels_295__flag;
	reg [0:0] ejection_channels_294__flag;
	reg [0:0] ejection_channels_293__flag;
	reg [0:0] ejection_channels_292__flag;
	reg [0:0] ejection_channels_291__flag;
	reg [0:0] ejection_channels_290__flag;
	reg [0:0] ejection_channels_289__flag;
	reg [0:0] ejection_channels_288__flag;
	reg [0:0] ejection_channels_287__flag;
	reg [0:0] ejection_channels_286__flag;
	reg [0:0] ejection_channels_285__flag;
	reg [0:0] ejection_channels_284__flag;
	reg [0:0] ejection_channels_283__flag;
	reg [0:0] ejection_channels_282__flag;
	reg [0:0] ejection_channels_281__flag;
	reg [0:0] ejection_channels_280__flag;
	reg [0:0] ejection_channels_279__flag;
	reg [0:0] ejection_channels_278__flag;
	reg [0:0] ejection_channels_277__flag;
	reg [0:0] ejection_channels_276__flag;
	reg [0:0] ejection_channels_275__flag;
	reg [0:0] ejection_channels_274__flag;
	reg [0:0] ejection_channels_273__flag;
	reg [0:0] ejection_channels_272__flag;
	reg [0:0] ejection_channels_271__flag;
	reg [0:0] ejection_channels_270__flag;
	reg [0:0] ejection_channels_269__flag;
	reg [0:0] ejection_channels_268__flag;
	reg [0:0] ejection_channels_267__flag;
	reg [0:0] ejection_channels_266__flag;
	reg [0:0] ejection_channels_265__flag;
	reg [0:0] ejection_channels_264__flag;
	reg [0:0] ejection_channels_263__flag;
	reg [0:0] ejection_channels_262__flag;
	reg [0:0] ejection_channels_261__flag;
	reg [0:0] ejection_channels_260__flag;
	reg [0:0] ejection_channels_259__flag;
	reg [0:0] ejection_channels_258__flag;
	reg [0:0] ejection_channels_257__flag;
	reg [0:0] ejection_channels_256__flag;
	reg [0:0] ejection_channels_255__flag;
	reg [0:0] ejection_channels_254__flag;
	reg [0:0] ejection_channels_253__flag;
	reg [0:0] ejection_channels_252__flag;
	reg [0:0] ejection_channels_251__flag;
	reg [0:0] ejection_channels_250__flag;
	reg [0:0] ejection_channels_249__flag;
	reg [0:0] ejection_channels_248__flag;
	reg [0:0] ejection_channels_247__flag;
	reg [0:0] ejection_channels_246__flag;
	reg [0:0] ejection_channels_245__flag;
	reg [0:0] ejection_channels_244__flag;
	reg [0:0] ejection_channels_243__flag;
	reg [0:0] ejection_channels_242__flag;
	reg [0:0] ejection_channels_241__flag;
	reg [0:0] ejection_channels_240__flag;
	reg [0:0] ejection_channels_239__flag;
	reg [0:0] ejection_channels_238__flag;
	reg [0:0] ejection_channels_237__flag;
	reg [0:0] ejection_channels_236__flag;
	reg [0:0] ejection_channels_235__flag;
	reg [0:0] ejection_channels_234__flag;
	reg [0:0] ejection_channels_233__flag;
	reg [0:0] ejection_channels_232__flag;
	reg [0:0] ejection_channels_231__flag;
	reg [0:0] ejection_channels_230__flag;
	reg [0:0] ejection_channels_229__flag;
	reg [0:0] ejection_channels_228__flag;
	reg [0:0] ejection_channels_227__flag;
	reg [0:0] ejection_channels_226__flag;
	reg [0:0] ejection_channels_225__flag;
	reg [0:0] ejection_channels_224__flag;
	reg [0:0] ejection_channels_223__flag;
	reg [0:0] ejection_channels_222__flag;
	reg [0:0] ejection_channels_221__flag;
	reg [0:0] ejection_channels_220__flag;
	reg [0:0] ejection_channels_219__flag;
	reg [0:0] ejection_channels_218__flag;
	reg [0:0] ejection_channels_217__flag;
	reg [0:0] ejection_channels_216__flag;
	reg [0:0] ejection_channels_215__flag;
	reg [0:0] ejection_channels_214__flag;
	reg [0:0] ejection_channels_213__flag;
	reg [0:0] ejection_channels_212__flag;
	reg [0:0] ejection_channels_211__flag;
	reg [0:0] ejection_channels_210__flag;
	reg [0:0] ejection_channels_209__flag;
	reg [0:0] ejection_channels_208__flag;
	reg [0:0] ejection_channels_207__flag;
	reg [0:0] ejection_channels_206__flag;
	reg [0:0] ejection_channels_205__flag;
	reg [0:0] ejection_channels_204__flag;
	reg [0:0] ejection_channels_203__flag;
	reg [0:0] ejection_channels_202__flag;
	reg [0:0] ejection_channels_201__flag;
	reg [0:0] ejection_channels_200__flag;
	reg [0:0] ejection_channels_199__flag;
	reg [0:0] ejection_channels_198__flag;
	reg [0:0] ejection_channels_197__flag;
	reg [0:0] ejection_channels_196__flag;
	reg [0:0] ejection_channels_195__flag;
	reg [0:0] ejection_channels_194__flag;
	reg [0:0] ejection_channels_193__flag;
	reg [0:0] ejection_channels_192__flag;
	reg [0:0] ejection_channels_191__flag;
	reg [0:0] ejection_channels_190__flag;
	reg [0:0] ejection_channels_189__flag;
	reg [0:0] ejection_channels_188__flag;
	reg [0:0] ejection_channels_187__flag;
	reg [0:0] ejection_channels_186__flag;
	reg [0:0] ejection_channels_185__flag;
	reg [0:0] ejection_channels_184__flag;
	reg [0:0] ejection_channels_183__flag;
	reg [0:0] ejection_channels_182__flag;
	reg [0:0] ejection_channels_181__flag;
	reg [0:0] ejection_channels_180__flag;
	reg [0:0] ejection_channels_179__flag;
	reg [0:0] ejection_channels_178__flag;
	reg [0:0] ejection_channels_177__flag;
	reg [0:0] ejection_channels_176__flag;
	reg [0:0] ejection_channels_175__flag;
	reg [0:0] ejection_channels_174__flag;
	reg [0:0] ejection_channels_173__flag;
	reg [0:0] ejection_channels_172__flag;
	reg [0:0] ejection_channels_171__flag;
	reg [0:0] ejection_channels_170__flag;
	reg [0:0] ejection_channels_169__flag;
	reg [0:0] ejection_channels_168__flag;
	reg [0:0] ejection_channels_167__flag;
	reg [0:0] ejection_channels_166__flag;
	reg [0:0] ejection_channels_165__flag;
	reg [0:0] ejection_channels_164__flag;
	reg [0:0] ejection_channels_163__flag;
	reg [0:0] ejection_channels_162__flag;
	reg [0:0] ejection_channels_161__flag;
	reg [0:0] ejection_channels_160__flag;
	reg [0:0] ejection_channels_159__flag;
	reg [0:0] ejection_channels_158__flag;
	reg [0:0] ejection_channels_157__flag;
	reg [0:0] ejection_channels_156__flag;
	reg [0:0] ejection_channels_155__flag;
	reg [0:0] ejection_channels_154__flag;
	reg [0:0] ejection_channels_153__flag;
	reg [0:0] ejection_channels_152__flag;
	reg [0:0] ejection_channels_151__flag;
	reg [0:0] ejection_channels_150__flag;
	reg [0:0] ejection_channels_149__flag;
	reg [0:0] ejection_channels_148__flag;
	reg [0:0] ejection_channels_147__flag;
	reg [0:0] ejection_channels_146__flag;
	reg [0:0] ejection_channels_145__flag;
	reg [0:0] ejection_channels_144__flag;
	reg [0:0] ejection_channels_143__flag;
	reg [0:0] ejection_channels_142__flag;
	reg [0:0] ejection_channels_141__flag;
	reg [0:0] ejection_channels_140__flag;
	reg [0:0] ejection_channels_139__flag;
	reg [0:0] ejection_channels_138__flag;
	reg [0:0] ejection_channels_137__flag;
	reg [0:0] ejection_channels_136__flag;
	reg [0:0] ejection_channels_135__flag;
	reg [0:0] ejection_channels_134__flag;
	reg [0:0] ejection_channels_133__flag;
	reg [0:0] ejection_channels_132__flag;
	reg [0:0] ejection_channels_131__flag;
	reg [0:0] ejection_channels_130__flag;
	reg [0:0] ejection_channels_129__flag;
	reg [0:0] ejection_channels_128__flag;
	reg [0:0] ejection_channels_127__flag;
	reg [0:0] ejection_channels_126__flag;
	reg [0:0] ejection_channels_125__flag;
	reg [0:0] ejection_channels_124__flag;
	reg [0:0] ejection_channels_123__flag;
	reg [0:0] ejection_channels_122__flag;
	reg [0:0] ejection_channels_121__flag;
	reg [0:0] ejection_channels_120__flag;
	reg [0:0] ejection_channels_119__flag;
	reg [0:0] ejection_channels_118__flag;
	reg [0:0] ejection_channels_117__flag;
	reg [0:0] ejection_channels_116__flag;
	reg [0:0] ejection_channels_115__flag;
	reg [0:0] ejection_channels_114__flag;
	reg [0:0] ejection_channels_113__flag;
	reg [0:0] ejection_channels_112__flag;
	reg [0:0] ejection_channels_111__flag;
	reg [0:0] ejection_channels_110__flag;
	reg [0:0] ejection_channels_109__flag;
	reg [0:0] ejection_channels_108__flag;
	reg [0:0] ejection_channels_107__flag;
	reg [0:0] ejection_channels_106__flag;
	reg [0:0] ejection_channels_105__flag;
	reg [0:0] ejection_channels_104__flag;
	reg [0:0] ejection_channels_103__flag;
	reg [0:0] ejection_channels_102__flag;
	reg [0:0] ejection_channels_101__flag;
	reg [0:0] ejection_channels_100__flag;
	reg [0:0] ejection_channels_99__flag;
	reg [0:0] ejection_channels_98__flag;
	reg [0:0] ejection_channels_97__flag;
	reg [0:0] ejection_channels_96__flag;
	reg [0:0] ejection_channels_95__flag;
	reg [0:0] ejection_channels_94__flag;
	reg [0:0] ejection_channels_93__flag;
	reg [0:0] ejection_channels_92__flag;
	reg [0:0] ejection_channels_91__flag;
	reg [0:0] ejection_channels_90__flag;
	reg [0:0] ejection_channels_89__flag;
	reg [0:0] ejection_channels_88__flag;
	reg [0:0] ejection_channels_87__flag;
	reg [0:0] ejection_channels_86__flag;
	reg [0:0] ejection_channels_85__flag;
	reg [0:0] ejection_channels_84__flag;
	reg [0:0] ejection_channels_83__flag;
	reg [0:0] ejection_channels_82__flag;
	reg [0:0] ejection_channels_81__flag;
	reg [0:0] ejection_channels_80__flag;
	reg [0:0] ejection_channels_79__flag;
	reg [0:0] ejection_channels_78__flag;
	reg [0:0] ejection_channels_77__flag;
	reg [0:0] ejection_channels_76__flag;
	reg [0:0] ejection_channels_75__flag;
	reg [0:0] ejection_channels_74__flag;
	reg [0:0] ejection_channels_73__flag;
	reg [0:0] ejection_channels_72__flag;
	reg [0:0] ejection_channels_71__flag;
	reg [0:0] ejection_channels_70__flag;
	reg [0:0] ejection_channels_69__flag;
	reg [0:0] ejection_channels_68__flag;
	reg [0:0] ejection_channels_67__flag;
	reg [0:0] ejection_channels_66__flag;
	reg [0:0] ejection_channels_65__flag;
	reg [0:0] ejection_channels_64__flag;
	reg [0:0] ejection_channels_63__flag;
	reg [0:0] ejection_channels_62__flag;
	reg [0:0] ejection_channels_61__flag;
	reg [0:0] ejection_channels_60__flag;
	reg [0:0] ejection_channels_59__flag;
	reg [0:0] ejection_channels_58__flag;
	reg [0:0] ejection_channels_57__flag;
	reg [0:0] ejection_channels_56__flag;
	reg [0:0] ejection_channels_55__flag;
	reg [0:0] ejection_channels_54__flag;
	reg [0:0] ejection_channels_53__flag;
	reg [0:0] ejection_channels_52__flag;
	reg [0:0] ejection_channels_51__flag;
	reg [0:0] ejection_channels_50__flag;
	reg [0:0] ejection_channels_49__flag;
	reg [0:0] ejection_channels_48__flag;
	reg [0:0] ejection_channels_47__flag;
	reg [0:0] ejection_channels_46__flag;
	reg [0:0] ejection_channels_45__flag;
	reg [0:0] ejection_channels_44__flag;
	reg [0:0] ejection_channels_43__flag;
	reg [0:0] ejection_channels_42__flag;
	reg [0:0] ejection_channels_41__flag;
	reg [0:0] ejection_channels_40__flag;
	reg [0:0] ejection_channels_39__flag;
	reg [0:0] ejection_channels_38__flag;
	reg [0:0] ejection_channels_37__flag;
	reg [0:0] ejection_channels_36__flag;
	reg [0:0] ejection_channels_35__flag;
	reg [0:0] ejection_channels_34__flag;
	reg [0:0] ejection_channels_33__flag;
	reg [0:0] ejection_channels_32__flag;
	reg [0:0] ejection_channels_31__flag;
	reg [0:0] ejection_channels_30__flag;
	reg [0:0] ejection_channels_29__flag;
	reg [0:0] ejection_channels_28__flag;
	reg [0:0] ejection_channels_27__flag;
	reg [0:0] ejection_channels_26__flag;
	reg [0:0] ejection_channels_25__flag;
	reg [0:0] ejection_channels_24__flag;
	reg [0:0] ejection_channels_23__flag;
	reg [0:0] ejection_channels_22__flag;
	reg [0:0] ejection_channels_21__flag;
	reg [0:0] ejection_channels_20__flag;
	reg [0:0] ejection_channels_19__flag;
	reg [0:0] ejection_channels_18__flag;
	reg [0:0] ejection_channels_17__flag;
	reg [0:0] ejection_channels_16__flag;
	reg [0:0] ejection_channels_15__flag;
	reg [0:0] ejection_channels_14__flag;
	reg [0:0] ejection_channels_13__flag;
	reg [0:0] ejection_channels_12__flag;
	reg [0:0] ejection_channels_11__flag;
	reg [0:0] ejection_channels_10__flag;
	reg [0:0] ejection_channels_9__flag;
	reg [0:0] ejection_channels_8__flag;
	reg [0:0] ejection_channels_7__flag;
	reg [0:0] ejection_channels_6__flag;
	reg [0:0] ejection_channels_5__flag;
	reg [0:0] ejection_channels_4__flag;
	reg [0:0] ejection_channels_3__flag;
	reg [0:0] ejection_channels_2__flag;
	reg [0:0] ejection_channels_1__flag;
	reg [0:0] ejection_channels_0__flag;
	reg [0:0] rtr_error_8__flag;
	reg [0:0] rtr_error_7__flag;
	reg [0:0] rtr_error_6__flag;
	reg [0:0] rtr_error_5__flag;
	reg [0:0] rtr_error_4__flag;
	reg [0:0] rtr_error_3__flag;
	reg [0:0] rtr_error_2__flag;
	reg [0:0] rtr_error_1__flag;
	reg [0:0] rtr_error_0__flag;

// ----- Error counter -------
	integer nb_error= 0;

// ----- FPGA fabric instanciation -------
	router_mesh_top_formal_verification FPGA_DUT(
		clk,
		reset,
		injection_channels_629_,
		injection_channels_628_,
		injection_channels_627_,
		injection_channels_626_,
		injection_channels_625_,
		injection_channels_624_,
		injection_channels_623_,
		injection_channels_622_,
		injection_channels_621_,
		injection_channels_620_,
		injection_channels_619_,
		injection_channels_618_,
		injection_channels_617_,
		injection_channels_616_,
		injection_channels_615_,
		injection_channels_614_,
		injection_channels_613_,
		injection_channels_612_,
		injection_channels_611_,
		injection_channels_610_,
		injection_channels_609_,
		injection_channels_608_,
		injection_channels_607_,
		injection_channels_606_,
		injection_channels_605_,
		injection_channels_604_,
		injection_channels_603_,
		injection_channels_602_,
		injection_channels_601_,
		injection_channels_600_,
		injection_channels_599_,
		injection_channels_598_,
		injection_channels_597_,
		injection_channels_596_,
		injection_channels_595_,
		injection_channels_594_,
		injection_channels_593_,
		injection_channels_592_,
		injection_channels_591_,
		injection_channels_590_,
		injection_channels_589_,
		injection_channels_588_,
		injection_channels_587_,
		injection_channels_586_,
		injection_channels_585_,
		injection_channels_584_,
		injection_channels_583_,
		injection_channels_582_,
		injection_channels_581_,
		injection_channels_580_,
		injection_channels_579_,
		injection_channels_578_,
		injection_channels_577_,
		injection_channels_576_,
		injection_channels_575_,
		injection_channels_574_,
		injection_channels_573_,
		injection_channels_572_,
		injection_channels_571_,
		injection_channels_570_,
		injection_channels_569_,
		injection_channels_568_,
		injection_channels_567_,
		injection_channels_566_,
		injection_channels_565_,
		injection_channels_564_,
		injection_channels_563_,
		injection_channels_562_,
		injection_channels_561_,
		injection_channels_560_,
		injection_channels_559_,
		injection_channels_558_,
		injection_channels_557_,
		injection_channels_556_,
		injection_channels_555_,
		injection_channels_554_,
		injection_channels_553_,
		injection_channels_552_,
		injection_channels_551_,
		injection_channels_550_,
		injection_channels_549_,
		injection_channels_548_,
		injection_channels_547_,
		injection_channels_546_,
		injection_channels_545_,
		injection_channels_544_,
		injection_channels_543_,
		injection_channels_542_,
		injection_channels_541_,
		injection_channels_540_,
		injection_channels_539_,
		injection_channels_538_,
		injection_channels_537_,
		injection_channels_536_,
		injection_channels_535_,
		injection_channels_534_,
		injection_channels_533_,
		injection_channels_532_,
		injection_channels_531_,
		injection_channels_530_,
		injection_channels_529_,
		injection_channels_528_,
		injection_channels_527_,
		injection_channels_526_,
		injection_channels_525_,
		injection_channels_524_,
		injection_channels_523_,
		injection_channels_522_,
		injection_channels_521_,
		injection_channels_520_,
		injection_channels_519_,
		injection_channels_518_,
		injection_channels_517_,
		injection_channels_516_,
		injection_channels_515_,
		injection_channels_514_,
		injection_channels_513_,
		injection_channels_512_,
		injection_channels_511_,
		injection_channels_510_,
		injection_channels_509_,
		injection_channels_508_,
		injection_channels_507_,
		injection_channels_506_,
		injection_channels_505_,
		injection_channels_504_,
		injection_channels_503_,
		injection_channels_502_,
		injection_channels_501_,
		injection_channels_500_,
		injection_channels_499_,
		injection_channels_498_,
		injection_channels_497_,
		injection_channels_496_,
		injection_channels_495_,
		injection_channels_494_,
		injection_channels_493_,
		injection_channels_492_,
		injection_channels_491_,
		injection_channels_490_,
		injection_channels_489_,
		injection_channels_488_,
		injection_channels_487_,
		injection_channels_486_,
		injection_channels_485_,
		injection_channels_484_,
		injection_channels_483_,
		injection_channels_482_,
		injection_channels_481_,
		injection_channels_480_,
		injection_channels_479_,
		injection_channels_478_,
		injection_channels_477_,
		injection_channels_476_,
		injection_channels_475_,
		injection_channels_474_,
		injection_channels_473_,
		injection_channels_472_,
		injection_channels_471_,
		injection_channels_470_,
		injection_channels_469_,
		injection_channels_468_,
		injection_channels_467_,
		injection_channels_466_,
		injection_channels_465_,
		injection_channels_464_,
		injection_channels_463_,
		injection_channels_462_,
		injection_channels_461_,
		injection_channels_460_,
		injection_channels_459_,
		injection_channels_458_,
		injection_channels_457_,
		injection_channels_456_,
		injection_channels_455_,
		injection_channels_454_,
		injection_channels_453_,
		injection_channels_452_,
		injection_channels_451_,
		injection_channels_450_,
		injection_channels_449_,
		injection_channels_448_,
		injection_channels_447_,
		injection_channels_446_,
		injection_channels_445_,
		injection_channels_444_,
		injection_channels_443_,
		injection_channels_442_,
		injection_channels_441_,
		injection_channels_440_,
		injection_channels_439_,
		injection_channels_438_,
		injection_channels_437_,
		injection_channels_436_,
		injection_channels_435_,
		injection_channels_434_,
		injection_channels_433_,
		injection_channels_432_,
		injection_channels_431_,
		injection_channels_430_,
		injection_channels_429_,
		injection_channels_428_,
		injection_channels_427_,
		injection_channels_426_,
		injection_channels_425_,
		injection_channels_424_,
		injection_channels_423_,
		injection_channels_422_,
		injection_channels_421_,
		injection_channels_420_,
		injection_channels_419_,
		injection_channels_418_,
		injection_channels_417_,
		injection_channels_416_,
		injection_channels_415_,
		injection_channels_414_,
		injection_channels_413_,
		injection_channels_412_,
		injection_channels_411_,
		injection_channels_410_,
		injection_channels_409_,
		injection_channels_408_,
		injection_channels_407_,
		injection_channels_406_,
		injection_channels_405_,
		injection_channels_404_,
		injection_channels_403_,
		injection_channels_402_,
		injection_channels_401_,
		injection_channels_400_,
		injection_channels_399_,
		injection_channels_398_,
		injection_channels_397_,
		injection_channels_396_,
		injection_channels_395_,
		injection_channels_394_,
		injection_channels_393_,
		injection_channels_392_,
		injection_channels_391_,
		injection_channels_390_,
		injection_channels_389_,
		injection_channels_388_,
		injection_channels_387_,
		injection_channels_386_,
		injection_channels_385_,
		injection_channels_384_,
		injection_channels_383_,
		injection_channels_382_,
		injection_channels_381_,
		injection_channels_380_,
		injection_channels_379_,
		injection_channels_378_,
		injection_channels_377_,
		injection_channels_376_,
		injection_channels_375_,
		injection_channels_374_,
		injection_channels_373_,
		injection_channels_372_,
		injection_channels_371_,
		injection_channels_370_,
		injection_channels_369_,
		injection_channels_368_,
		injection_channels_367_,
		injection_channels_366_,
		injection_channels_365_,
		injection_channels_364_,
		injection_channels_363_,
		injection_channels_362_,
		injection_channels_361_,
		injection_channels_360_,
		injection_channels_359_,
		injection_channels_358_,
		injection_channels_357_,
		injection_channels_356_,
		injection_channels_355_,
		injection_channels_354_,
		injection_channels_353_,
		injection_channels_352_,
		injection_channels_351_,
		injection_channels_350_,
		injection_channels_349_,
		injection_channels_348_,
		injection_channels_347_,
		injection_channels_346_,
		injection_channels_345_,
		injection_channels_344_,
		injection_channels_343_,
		injection_channels_342_,
		injection_channels_341_,
		injection_channels_340_,
		injection_channels_339_,
		injection_channels_338_,
		injection_channels_337_,
		injection_channels_336_,
		injection_channels_335_,
		injection_channels_334_,
		injection_channels_333_,
		injection_channels_332_,
		injection_channels_331_,
		injection_channels_330_,
		injection_channels_329_,
		injection_channels_328_,
		injection_channels_327_,
		injection_channels_326_,
		injection_channels_325_,
		injection_channels_324_,
		injection_channels_323_,
		injection_channels_322_,
		injection_channels_321_,
		injection_channels_320_,
		injection_channels_319_,
		injection_channels_318_,
		injection_channels_317_,
		injection_channels_316_,
		injection_channels_315_,
		injection_channels_314_,
		injection_channels_313_,
		injection_channels_312_,
		injection_channels_311_,
		injection_channels_310_,
		injection_channels_309_,
		injection_channels_308_,
		injection_channels_307_,
		injection_channels_306_,
		injection_channels_305_,
		injection_channels_304_,
		injection_channels_303_,
		injection_channels_302_,
		injection_channels_301_,
		injection_channels_300_,
		injection_channels_299_,
		injection_channels_298_,
		injection_channels_297_,
		injection_channels_296_,
		injection_channels_295_,
		injection_channels_294_,
		injection_channels_293_,
		injection_channels_292_,
		injection_channels_291_,
		injection_channels_290_,
		injection_channels_289_,
		injection_channels_288_,
		injection_channels_287_,
		injection_channels_286_,
		injection_channels_285_,
		injection_channels_284_,
		injection_channels_283_,
		injection_channels_282_,
		injection_channels_281_,
		injection_channels_280_,
		injection_channels_279_,
		injection_channels_278_,
		injection_channels_277_,
		injection_channels_276_,
		injection_channels_275_,
		injection_channels_274_,
		injection_channels_273_,
		injection_channels_272_,
		injection_channels_271_,
		injection_channels_270_,
		injection_channels_269_,
		injection_channels_268_,
		injection_channels_267_,
		injection_channels_266_,
		injection_channels_265_,
		injection_channels_264_,
		injection_channels_263_,
		injection_channels_262_,
		injection_channels_261_,
		injection_channels_260_,
		injection_channels_259_,
		injection_channels_258_,
		injection_channels_257_,
		injection_channels_256_,
		injection_channels_255_,
		injection_channels_254_,
		injection_channels_253_,
		injection_channels_252_,
		injection_channels_251_,
		injection_channels_250_,
		injection_channels_249_,
		injection_channels_248_,
		injection_channels_247_,
		injection_channels_246_,
		injection_channels_245_,
		injection_channels_244_,
		injection_channels_243_,
		injection_channels_242_,
		injection_channels_241_,
		injection_channels_240_,
		injection_channels_239_,
		injection_channels_238_,
		injection_channels_237_,
		injection_channels_236_,
		injection_channels_235_,
		injection_channels_234_,
		injection_channels_233_,
		injection_channels_232_,
		injection_channels_231_,
		injection_channels_230_,
		injection_channels_229_,
		injection_channels_228_,
		injection_channels_227_,
		injection_channels_226_,
		injection_channels_225_,
		injection_channels_224_,
		injection_channels_223_,
		injection_channels_222_,
		injection_channels_221_,
		injection_channels_220_,
		injection_channels_219_,
		injection_channels_218_,
		injection_channels_217_,
		injection_channels_216_,
		injection_channels_215_,
		injection_channels_214_,
		injection_channels_213_,
		injection_channels_212_,
		injection_channels_211_,
		injection_channels_210_,
		injection_channels_209_,
		injection_channels_208_,
		injection_channels_207_,
		injection_channels_206_,
		injection_channels_205_,
		injection_channels_204_,
		injection_channels_203_,
		injection_channels_202_,
		injection_channels_201_,
		injection_channels_200_,
		injection_channels_199_,
		injection_channels_198_,
		injection_channels_197_,
		injection_channels_196_,
		injection_channels_195_,
		injection_channels_194_,
		injection_channels_193_,
		injection_channels_192_,
		injection_channels_191_,
		injection_channels_190_,
		injection_channels_189_,
		injection_channels_188_,
		injection_channels_187_,
		injection_channels_186_,
		injection_channels_185_,
		injection_channels_184_,
		injection_channels_183_,
		injection_channels_182_,
		injection_channels_181_,
		injection_channels_180_,
		injection_channels_179_,
		injection_channels_178_,
		injection_channels_177_,
		injection_channels_176_,
		injection_channels_175_,
		injection_channels_174_,
		injection_channels_173_,
		injection_channels_172_,
		injection_channels_171_,
		injection_channels_170_,
		injection_channels_169_,
		injection_channels_168_,
		injection_channels_167_,
		injection_channels_166_,
		injection_channels_165_,
		injection_channels_164_,
		injection_channels_163_,
		injection_channels_162_,
		injection_channels_161_,
		injection_channels_160_,
		injection_channels_159_,
		injection_channels_158_,
		injection_channels_157_,
		injection_channels_156_,
		injection_channels_155_,
		injection_channels_154_,
		injection_channels_153_,
		injection_channels_152_,
		injection_channels_151_,
		injection_channels_150_,
		injection_channels_149_,
		injection_channels_148_,
		injection_channels_147_,
		injection_channels_146_,
		injection_channels_145_,
		injection_channels_144_,
		injection_channels_143_,
		injection_channels_142_,
		injection_channels_141_,
		injection_channels_140_,
		injection_channels_139_,
		injection_channels_138_,
		injection_channels_137_,
		injection_channels_136_,
		injection_channels_135_,
		injection_channels_134_,
		injection_channels_133_,
		injection_channels_132_,
		injection_channels_131_,
		injection_channels_130_,
		injection_channels_129_,
		injection_channels_128_,
		injection_channels_127_,
		injection_channels_126_,
		injection_channels_125_,
		injection_channels_124_,
		injection_channels_123_,
		injection_channels_122_,
		injection_channels_121_,
		injection_channels_120_,
		injection_channels_119_,
		injection_channels_118_,
		injection_channels_117_,
		injection_channels_116_,
		injection_channels_115_,
		injection_channels_114_,
		injection_channels_113_,
		injection_channels_112_,
		injection_channels_111_,
		injection_channels_110_,
		injection_channels_109_,
		injection_channels_108_,
		injection_channels_107_,
		injection_channels_106_,
		injection_channels_105_,
		injection_channels_104_,
		injection_channels_103_,
		injection_channels_102_,
		injection_channels_101_,
		injection_channels_100_,
		injection_channels_99_,
		injection_channels_98_,
		injection_channels_97_,
		injection_channels_96_,
		injection_channels_95_,
		injection_channels_94_,
		injection_channels_93_,
		injection_channels_92_,
		injection_channels_91_,
		injection_channels_90_,
		injection_channels_89_,
		injection_channels_88_,
		injection_channels_87_,
		injection_channels_86_,
		injection_channels_85_,
		injection_channels_84_,
		injection_channels_83_,
		injection_channels_82_,
		injection_channels_81_,
		injection_channels_80_,
		injection_channels_79_,
		injection_channels_78_,
		injection_channels_77_,
		injection_channels_76_,
		injection_channels_75_,
		injection_channels_74_,
		injection_channels_73_,
		injection_channels_72_,
		injection_channels_71_,
		injection_channels_70_,
		injection_channels_69_,
		injection_channels_68_,
		injection_channels_67_,
		injection_channels_66_,
		injection_channels_65_,
		injection_channels_64_,
		injection_channels_63_,
		injection_channels_62_,
		injection_channels_61_,
		injection_channels_60_,
		injection_channels_59_,
		injection_channels_58_,
		injection_channels_57_,
		injection_channels_56_,
		injection_channels_55_,
		injection_channels_54_,
		injection_channels_53_,
		injection_channels_52_,
		injection_channels_51_,
		injection_channels_50_,
		injection_channels_49_,
		injection_channels_48_,
		injection_channels_47_,
		injection_channels_46_,
		injection_channels_45_,
		injection_channels_44_,
		injection_channels_43_,
		injection_channels_42_,
		injection_channels_41_,
		injection_channels_40_,
		injection_channels_39_,
		injection_channels_38_,
		injection_channels_37_,
		injection_channels_36_,
		injection_channels_35_,
		injection_channels_34_,
		injection_channels_33_,
		injection_channels_32_,
		injection_channels_31_,
		injection_channels_30_,
		injection_channels_29_,
		injection_channels_28_,
		injection_channels_27_,
		injection_channels_26_,
		injection_channels_25_,
		injection_channels_24_,
		injection_channels_23_,
		injection_channels_22_,
		injection_channels_21_,
		injection_channels_20_,
		injection_channels_19_,
		injection_channels_18_,
		injection_channels_17_,
		injection_channels_16_,
		injection_channels_15_,
		injection_channels_14_,
		injection_channels_13_,
		injection_channels_12_,
		injection_channels_11_,
		injection_channels_10_,
		injection_channels_9_,
		injection_channels_8_,
		injection_channels_7_,
		injection_channels_6_,
		injection_channels_5_,
		injection_channels_4_,
		injection_channels_3_,
		injection_channels_2_,
		injection_channels_1_,
		injection_channels_0_,
		ejection_flow_ctrl_26_,
		ejection_flow_ctrl_25_,
		ejection_flow_ctrl_24_,
		ejection_flow_ctrl_23_,
		ejection_flow_ctrl_22_,
		ejection_flow_ctrl_21_,
		ejection_flow_ctrl_20_,
		ejection_flow_ctrl_19_,
		ejection_flow_ctrl_18_,
		ejection_flow_ctrl_17_,
		ejection_flow_ctrl_16_,
		ejection_flow_ctrl_15_,
		ejection_flow_ctrl_14_,
		ejection_flow_ctrl_13_,
		ejection_flow_ctrl_12_,
		ejection_flow_ctrl_11_,
		ejection_flow_ctrl_10_,
		ejection_flow_ctrl_9_,
		ejection_flow_ctrl_8_,
		ejection_flow_ctrl_7_,
		ejection_flow_ctrl_6_,
		ejection_flow_ctrl_5_,
		ejection_flow_ctrl_4_,
		ejection_flow_ctrl_3_,
		ejection_flow_ctrl_2_,
		ejection_flow_ctrl_1_,
		ejection_flow_ctrl_0_,
		injection_flow_ctrl_26__gfpga,
		injection_flow_ctrl_25__gfpga,
		injection_flow_ctrl_24__gfpga,
		injection_flow_ctrl_23__gfpga,
		injection_flow_ctrl_22__gfpga,
		injection_flow_ctrl_21__gfpga,
		injection_flow_ctrl_20__gfpga,
		injection_flow_ctrl_19__gfpga,
		injection_flow_ctrl_18__gfpga,
		injection_flow_ctrl_17__gfpga,
		injection_flow_ctrl_16__gfpga,
		injection_flow_ctrl_15__gfpga,
		injection_flow_ctrl_14__gfpga,
		injection_flow_ctrl_13__gfpga,
		injection_flow_ctrl_12__gfpga,
		injection_flow_ctrl_11__gfpga,
		injection_flow_ctrl_10__gfpga,
		injection_flow_ctrl_9__gfpga,
		injection_flow_ctrl_8__gfpga,
		injection_flow_ctrl_7__gfpga,
		injection_flow_ctrl_6__gfpga,
		injection_flow_ctrl_5__gfpga,
		injection_flow_ctrl_4__gfpga,
		injection_flow_ctrl_3__gfpga,
		injection_flow_ctrl_2__gfpga,
		injection_flow_ctrl_1__gfpga,
		injection_flow_ctrl_0__gfpga,
		ejection_channels_629__gfpga,
		ejection_channels_628__gfpga,
		ejection_channels_627__gfpga,
		ejection_channels_626__gfpga,
		ejection_channels_625__gfpga,
		ejection_channels_624__gfpga,
		ejection_channels_623__gfpga,
		ejection_channels_622__gfpga,
		ejection_channels_621__gfpga,
		ejection_channels_620__gfpga,
		ejection_channels_619__gfpga,
		ejection_channels_618__gfpga,
		ejection_channels_617__gfpga,
		ejection_channels_616__gfpga,
		ejection_channels_615__gfpga,
		ejection_channels_614__gfpga,
		ejection_channels_613__gfpga,
		ejection_channels_612__gfpga,
		ejection_channels_611__gfpga,
		ejection_channels_610__gfpga,
		ejection_channels_609__gfpga,
		ejection_channels_608__gfpga,
		ejection_channels_607__gfpga,
		ejection_channels_606__gfpga,
		ejection_channels_605__gfpga,
		ejection_channels_604__gfpga,
		ejection_channels_603__gfpga,
		ejection_channels_602__gfpga,
		ejection_channels_601__gfpga,
		ejection_channels_600__gfpga,
		ejection_channels_599__gfpga,
		ejection_channels_598__gfpga,
		ejection_channels_597__gfpga,
		ejection_channels_596__gfpga,
		ejection_channels_595__gfpga,
		ejection_channels_594__gfpga,
		ejection_channels_593__gfpga,
		ejection_channels_592__gfpga,
		ejection_channels_591__gfpga,
		ejection_channels_590__gfpga,
		ejection_channels_589__gfpga,
		ejection_channels_588__gfpga,
		ejection_channels_587__gfpga,
		ejection_channels_586__gfpga,
		ejection_channels_585__gfpga,
		ejection_channels_584__gfpga,
		ejection_channels_583__gfpga,
		ejection_channels_582__gfpga,
		ejection_channels_581__gfpga,
		ejection_channels_580__gfpga,
		ejection_channels_579__gfpga,
		ejection_channels_578__gfpga,
		ejection_channels_577__gfpga,
		ejection_channels_576__gfpga,
		ejection_channels_575__gfpga,
		ejection_channels_574__gfpga,
		ejection_channels_573__gfpga,
		ejection_channels_572__gfpga,
		ejection_channels_571__gfpga,
		ejection_channels_570__gfpga,
		ejection_channels_569__gfpga,
		ejection_channels_568__gfpga,
		ejection_channels_567__gfpga,
		ejection_channels_566__gfpga,
		ejection_channels_565__gfpga,
		ejection_channels_564__gfpga,
		ejection_channels_563__gfpga,
		ejection_channels_562__gfpga,
		ejection_channels_561__gfpga,
		ejection_channels_560__gfpga,
		ejection_channels_559__gfpga,
		ejection_channels_558__gfpga,
		ejection_channels_557__gfpga,
		ejection_channels_556__gfpga,
		ejection_channels_555__gfpga,
		ejection_channels_554__gfpga,
		ejection_channels_553__gfpga,
		ejection_channels_552__gfpga,
		ejection_channels_551__gfpga,
		ejection_channels_550__gfpga,
		ejection_channels_549__gfpga,
		ejection_channels_548__gfpga,
		ejection_channels_547__gfpga,
		ejection_channels_546__gfpga,
		ejection_channels_545__gfpga,
		ejection_channels_544__gfpga,
		ejection_channels_543__gfpga,
		ejection_channels_542__gfpga,
		ejection_channels_541__gfpga,
		ejection_channels_540__gfpga,
		ejection_channels_539__gfpga,
		ejection_channels_538__gfpga,
		ejection_channels_537__gfpga,
		ejection_channels_536__gfpga,
		ejection_channels_535__gfpga,
		ejection_channels_534__gfpga,
		ejection_channels_533__gfpga,
		ejection_channels_532__gfpga,
		ejection_channels_531__gfpga,
		ejection_channels_530__gfpga,
		ejection_channels_529__gfpga,
		ejection_channels_528__gfpga,
		ejection_channels_527__gfpga,
		ejection_channels_526__gfpga,
		ejection_channels_525__gfpga,
		ejection_channels_524__gfpga,
		ejection_channels_523__gfpga,
		ejection_channels_522__gfpga,
		ejection_channels_521__gfpga,
		ejection_channels_520__gfpga,
		ejection_channels_519__gfpga,
		ejection_channels_518__gfpga,
		ejection_channels_517__gfpga,
		ejection_channels_516__gfpga,
		ejection_channels_515__gfpga,
		ejection_channels_514__gfpga,
		ejection_channels_513__gfpga,
		ejection_channels_512__gfpga,
		ejection_channels_511__gfpga,
		ejection_channels_510__gfpga,
		ejection_channels_509__gfpga,
		ejection_channels_508__gfpga,
		ejection_channels_507__gfpga,
		ejection_channels_506__gfpga,
		ejection_channels_505__gfpga,
		ejection_channels_504__gfpga,
		ejection_channels_503__gfpga,
		ejection_channels_502__gfpga,
		ejection_channels_501__gfpga,
		ejection_channels_500__gfpga,
		ejection_channels_499__gfpga,
		ejection_channels_498__gfpga,
		ejection_channels_497__gfpga,
		ejection_channels_496__gfpga,
		ejection_channels_495__gfpga,
		ejection_channels_494__gfpga,
		ejection_channels_493__gfpga,
		ejection_channels_492__gfpga,
		ejection_channels_491__gfpga,
		ejection_channels_490__gfpga,
		ejection_channels_489__gfpga,
		ejection_channels_488__gfpga,
		ejection_channels_487__gfpga,
		ejection_channels_486__gfpga,
		ejection_channels_485__gfpga,
		ejection_channels_484__gfpga,
		ejection_channels_483__gfpga,
		ejection_channels_482__gfpga,
		ejection_channels_481__gfpga,
		ejection_channels_480__gfpga,
		ejection_channels_479__gfpga,
		ejection_channels_478__gfpga,
		ejection_channels_477__gfpga,
		ejection_channels_476__gfpga,
		ejection_channels_475__gfpga,
		ejection_channels_474__gfpga,
		ejection_channels_473__gfpga,
		ejection_channels_472__gfpga,
		ejection_channels_471__gfpga,
		ejection_channels_470__gfpga,
		ejection_channels_469__gfpga,
		ejection_channels_468__gfpga,
		ejection_channels_467__gfpga,
		ejection_channels_466__gfpga,
		ejection_channels_465__gfpga,
		ejection_channels_464__gfpga,
		ejection_channels_463__gfpga,
		ejection_channels_462__gfpga,
		ejection_channels_461__gfpga,
		ejection_channels_460__gfpga,
		ejection_channels_459__gfpga,
		ejection_channels_458__gfpga,
		ejection_channels_457__gfpga,
		ejection_channels_456__gfpga,
		ejection_channels_455__gfpga,
		ejection_channels_454__gfpga,
		ejection_channels_453__gfpga,
		ejection_channels_452__gfpga,
		ejection_channels_451__gfpga,
		ejection_channels_450__gfpga,
		ejection_channels_449__gfpga,
		ejection_channels_448__gfpga,
		ejection_channels_447__gfpga,
		ejection_channels_446__gfpga,
		ejection_channels_445__gfpga,
		ejection_channels_444__gfpga,
		ejection_channels_443__gfpga,
		ejection_channels_442__gfpga,
		ejection_channels_441__gfpga,
		ejection_channels_440__gfpga,
		ejection_channels_439__gfpga,
		ejection_channels_438__gfpga,
		ejection_channels_437__gfpga,
		ejection_channels_436__gfpga,
		ejection_channels_435__gfpga,
		ejection_channels_434__gfpga,
		ejection_channels_433__gfpga,
		ejection_channels_432__gfpga,
		ejection_channels_431__gfpga,
		ejection_channels_430__gfpga,
		ejection_channels_429__gfpga,
		ejection_channels_428__gfpga,
		ejection_channels_427__gfpga,
		ejection_channels_426__gfpga,
		ejection_channels_425__gfpga,
		ejection_channels_424__gfpga,
		ejection_channels_423__gfpga,
		ejection_channels_422__gfpga,
		ejection_channels_421__gfpga,
		ejection_channels_420__gfpga,
		ejection_channels_419__gfpga,
		ejection_channels_418__gfpga,
		ejection_channels_417__gfpga,
		ejection_channels_416__gfpga,
		ejection_channels_415__gfpga,
		ejection_channels_414__gfpga,
		ejection_channels_413__gfpga,
		ejection_channels_412__gfpga,
		ejection_channels_411__gfpga,
		ejection_channels_410__gfpga,
		ejection_channels_409__gfpga,
		ejection_channels_408__gfpga,
		ejection_channels_407__gfpga,
		ejection_channels_406__gfpga,
		ejection_channels_405__gfpga,
		ejection_channels_404__gfpga,
		ejection_channels_403__gfpga,
		ejection_channels_402__gfpga,
		ejection_channels_401__gfpga,
		ejection_channels_400__gfpga,
		ejection_channels_399__gfpga,
		ejection_channels_398__gfpga,
		ejection_channels_397__gfpga,
		ejection_channels_396__gfpga,
		ejection_channels_395__gfpga,
		ejection_channels_394__gfpga,
		ejection_channels_393__gfpga,
		ejection_channels_392__gfpga,
		ejection_channels_391__gfpga,
		ejection_channels_390__gfpga,
		ejection_channels_389__gfpga,
		ejection_channels_388__gfpga,
		ejection_channels_387__gfpga,
		ejection_channels_386__gfpga,
		ejection_channels_385__gfpga,
		ejection_channels_384__gfpga,
		ejection_channels_383__gfpga,
		ejection_channels_382__gfpga,
		ejection_channels_381__gfpga,
		ejection_channels_380__gfpga,
		ejection_channels_379__gfpga,
		ejection_channels_378__gfpga,
		ejection_channels_377__gfpga,
		ejection_channels_376__gfpga,
		ejection_channels_375__gfpga,
		ejection_channels_374__gfpga,
		ejection_channels_373__gfpga,
		ejection_channels_372__gfpga,
		ejection_channels_371__gfpga,
		ejection_channels_370__gfpga,
		ejection_channels_369__gfpga,
		ejection_channels_368__gfpga,
		ejection_channels_367__gfpga,
		ejection_channels_366__gfpga,
		ejection_channels_365__gfpga,
		ejection_channels_364__gfpga,
		ejection_channels_363__gfpga,
		ejection_channels_362__gfpga,
		ejection_channels_361__gfpga,
		ejection_channels_360__gfpga,
		ejection_channels_359__gfpga,
		ejection_channels_358__gfpga,
		ejection_channels_357__gfpga,
		ejection_channels_356__gfpga,
		ejection_channels_355__gfpga,
		ejection_channels_354__gfpga,
		ejection_channels_353__gfpga,
		ejection_channels_352__gfpga,
		ejection_channels_351__gfpga,
		ejection_channels_350__gfpga,
		ejection_channels_349__gfpga,
		ejection_channels_348__gfpga,
		ejection_channels_347__gfpga,
		ejection_channels_346__gfpga,
		ejection_channels_345__gfpga,
		ejection_channels_344__gfpga,
		ejection_channels_343__gfpga,
		ejection_channels_342__gfpga,
		ejection_channels_341__gfpga,
		ejection_channels_340__gfpga,
		ejection_channels_339__gfpga,
		ejection_channels_338__gfpga,
		ejection_channels_337__gfpga,
		ejection_channels_336__gfpga,
		ejection_channels_335__gfpga,
		ejection_channels_334__gfpga,
		ejection_channels_333__gfpga,
		ejection_channels_332__gfpga,
		ejection_channels_331__gfpga,
		ejection_channels_330__gfpga,
		ejection_channels_329__gfpga,
		ejection_channels_328__gfpga,
		ejection_channels_327__gfpga,
		ejection_channels_326__gfpga,
		ejection_channels_325__gfpga,
		ejection_channels_324__gfpga,
		ejection_channels_323__gfpga,
		ejection_channels_322__gfpga,
		ejection_channels_321__gfpga,
		ejection_channels_320__gfpga,
		ejection_channels_319__gfpga,
		ejection_channels_318__gfpga,
		ejection_channels_317__gfpga,
		ejection_channels_316__gfpga,
		ejection_channels_315__gfpga,
		ejection_channels_314__gfpga,
		ejection_channels_313__gfpga,
		ejection_channels_312__gfpga,
		ejection_channels_311__gfpga,
		ejection_channels_310__gfpga,
		ejection_channels_309__gfpga,
		ejection_channels_308__gfpga,
		ejection_channels_307__gfpga,
		ejection_channels_306__gfpga,
		ejection_channels_305__gfpga,
		ejection_channels_304__gfpga,
		ejection_channels_303__gfpga,
		ejection_channels_302__gfpga,
		ejection_channels_301__gfpga,
		ejection_channels_300__gfpga,
		ejection_channels_299__gfpga,
		ejection_channels_298__gfpga,
		ejection_channels_297__gfpga,
		ejection_channels_296__gfpga,
		ejection_channels_295__gfpga,
		ejection_channels_294__gfpga,
		ejection_channels_293__gfpga,
		ejection_channels_292__gfpga,
		ejection_channels_291__gfpga,
		ejection_channels_290__gfpga,
		ejection_channels_289__gfpga,
		ejection_channels_288__gfpga,
		ejection_channels_287__gfpga,
		ejection_channels_286__gfpga,
		ejection_channels_285__gfpga,
		ejection_channels_284__gfpga,
		ejection_channels_283__gfpga,
		ejection_channels_282__gfpga,
		ejection_channels_281__gfpga,
		ejection_channels_280__gfpga,
		ejection_channels_279__gfpga,
		ejection_channels_278__gfpga,
		ejection_channels_277__gfpga,
		ejection_channels_276__gfpga,
		ejection_channels_275__gfpga,
		ejection_channels_274__gfpga,
		ejection_channels_273__gfpga,
		ejection_channels_272__gfpga,
		ejection_channels_271__gfpga,
		ejection_channels_270__gfpga,
		ejection_channels_269__gfpga,
		ejection_channels_268__gfpga,
		ejection_channels_267__gfpga,
		ejection_channels_266__gfpga,
		ejection_channels_265__gfpga,
		ejection_channels_264__gfpga,
		ejection_channels_263__gfpga,
		ejection_channels_262__gfpga,
		ejection_channels_261__gfpga,
		ejection_channels_260__gfpga,
		ejection_channels_259__gfpga,
		ejection_channels_258__gfpga,
		ejection_channels_257__gfpga,
		ejection_channels_256__gfpga,
		ejection_channels_255__gfpga,
		ejection_channels_254__gfpga,
		ejection_channels_253__gfpga,
		ejection_channels_252__gfpga,
		ejection_channels_251__gfpga,
		ejection_channels_250__gfpga,
		ejection_channels_249__gfpga,
		ejection_channels_248__gfpga,
		ejection_channels_247__gfpga,
		ejection_channels_246__gfpga,
		ejection_channels_245__gfpga,
		ejection_channels_244__gfpga,
		ejection_channels_243__gfpga,
		ejection_channels_242__gfpga,
		ejection_channels_241__gfpga,
		ejection_channels_240__gfpga,
		ejection_channels_239__gfpga,
		ejection_channels_238__gfpga,
		ejection_channels_237__gfpga,
		ejection_channels_236__gfpga,
		ejection_channels_235__gfpga,
		ejection_channels_234__gfpga,
		ejection_channels_233__gfpga,
		ejection_channels_232__gfpga,
		ejection_channels_231__gfpga,
		ejection_channels_230__gfpga,
		ejection_channels_229__gfpga,
		ejection_channels_228__gfpga,
		ejection_channels_227__gfpga,
		ejection_channels_226__gfpga,
		ejection_channels_225__gfpga,
		ejection_channels_224__gfpga,
		ejection_channels_223__gfpga,
		ejection_channels_222__gfpga,
		ejection_channels_221__gfpga,
		ejection_channels_220__gfpga,
		ejection_channels_219__gfpga,
		ejection_channels_218__gfpga,
		ejection_channels_217__gfpga,
		ejection_channels_216__gfpga,
		ejection_channels_215__gfpga,
		ejection_channels_214__gfpga,
		ejection_channels_213__gfpga,
		ejection_channels_212__gfpga,
		ejection_channels_211__gfpga,
		ejection_channels_210__gfpga,
		ejection_channels_209__gfpga,
		ejection_channels_208__gfpga,
		ejection_channels_207__gfpga,
		ejection_channels_206__gfpga,
		ejection_channels_205__gfpga,
		ejection_channels_204__gfpga,
		ejection_channels_203__gfpga,
		ejection_channels_202__gfpga,
		ejection_channels_201__gfpga,
		ejection_channels_200__gfpga,
		ejection_channels_199__gfpga,
		ejection_channels_198__gfpga,
		ejection_channels_197__gfpga,
		ejection_channels_196__gfpga,
		ejection_channels_195__gfpga,
		ejection_channels_194__gfpga,
		ejection_channels_193__gfpga,
		ejection_channels_192__gfpga,
		ejection_channels_191__gfpga,
		ejection_channels_190__gfpga,
		ejection_channels_189__gfpga,
		ejection_channels_188__gfpga,
		ejection_channels_187__gfpga,
		ejection_channels_186__gfpga,
		ejection_channels_185__gfpga,
		ejection_channels_184__gfpga,
		ejection_channels_183__gfpga,
		ejection_channels_182__gfpga,
		ejection_channels_181__gfpga,
		ejection_channels_180__gfpga,
		ejection_channels_179__gfpga,
		ejection_channels_178__gfpga,
		ejection_channels_177__gfpga,
		ejection_channels_176__gfpga,
		ejection_channels_175__gfpga,
		ejection_channels_174__gfpga,
		ejection_channels_173__gfpga,
		ejection_channels_172__gfpga,
		ejection_channels_171__gfpga,
		ejection_channels_170__gfpga,
		ejection_channels_169__gfpga,
		ejection_channels_168__gfpga,
		ejection_channels_167__gfpga,
		ejection_channels_166__gfpga,
		ejection_channels_165__gfpga,
		ejection_channels_164__gfpga,
		ejection_channels_163__gfpga,
		ejection_channels_162__gfpga,
		ejection_channels_161__gfpga,
		ejection_channels_160__gfpga,
		ejection_channels_159__gfpga,
		ejection_channels_158__gfpga,
		ejection_channels_157__gfpga,
		ejection_channels_156__gfpga,
		ejection_channels_155__gfpga,
		ejection_channels_154__gfpga,
		ejection_channels_153__gfpga,
		ejection_channels_152__gfpga,
		ejection_channels_151__gfpga,
		ejection_channels_150__gfpga,
		ejection_channels_149__gfpga,
		ejection_channels_148__gfpga,
		ejection_channels_147__gfpga,
		ejection_channels_146__gfpga,
		ejection_channels_145__gfpga,
		ejection_channels_144__gfpga,
		ejection_channels_143__gfpga,
		ejection_channels_142__gfpga,
		ejection_channels_141__gfpga,
		ejection_channels_140__gfpga,
		ejection_channels_139__gfpga,
		ejection_channels_138__gfpga,
		ejection_channels_137__gfpga,
		ejection_channels_136__gfpga,
		ejection_channels_135__gfpga,
		ejection_channels_134__gfpga,
		ejection_channels_133__gfpga,
		ejection_channels_132__gfpga,
		ejection_channels_131__gfpga,
		ejection_channels_130__gfpga,
		ejection_channels_129__gfpga,
		ejection_channels_128__gfpga,
		ejection_channels_127__gfpga,
		ejection_channels_126__gfpga,
		ejection_channels_125__gfpga,
		ejection_channels_124__gfpga,
		ejection_channels_123__gfpga,
		ejection_channels_122__gfpga,
		ejection_channels_121__gfpga,
		ejection_channels_120__gfpga,
		ejection_channels_119__gfpga,
		ejection_channels_118__gfpga,
		ejection_channels_117__gfpga,
		ejection_channels_116__gfpga,
		ejection_channels_115__gfpga,
		ejection_channels_114__gfpga,
		ejection_channels_113__gfpga,
		ejection_channels_112__gfpga,
		ejection_channels_111__gfpga,
		ejection_channels_110__gfpga,
		ejection_channels_109__gfpga,
		ejection_channels_108__gfpga,
		ejection_channels_107__gfpga,
		ejection_channels_106__gfpga,
		ejection_channels_105__gfpga,
		ejection_channels_104__gfpga,
		ejection_channels_103__gfpga,
		ejection_channels_102__gfpga,
		ejection_channels_101__gfpga,
		ejection_channels_100__gfpga,
		ejection_channels_99__gfpga,
		ejection_channels_98__gfpga,
		ejection_channels_97__gfpga,
		ejection_channels_96__gfpga,
		ejection_channels_95__gfpga,
		ejection_channels_94__gfpga,
		ejection_channels_93__gfpga,
		ejection_channels_92__gfpga,
		ejection_channels_91__gfpga,
		ejection_channels_90__gfpga,
		ejection_channels_89__gfpga,
		ejection_channels_88__gfpga,
		ejection_channels_87__gfpga,
		ejection_channels_86__gfpga,
		ejection_channels_85__gfpga,
		ejection_channels_84__gfpga,
		ejection_channels_83__gfpga,
		ejection_channels_82__gfpga,
		ejection_channels_81__gfpga,
		ejection_channels_80__gfpga,
		ejection_channels_79__gfpga,
		ejection_channels_78__gfpga,
		ejection_channels_77__gfpga,
		ejection_channels_76__gfpga,
		ejection_channels_75__gfpga,
		ejection_channels_74__gfpga,
		ejection_channels_73__gfpga,
		ejection_channels_72__gfpga,
		ejection_channels_71__gfpga,
		ejection_channels_70__gfpga,
		ejection_channels_69__gfpga,
		ejection_channels_68__gfpga,
		ejection_channels_67__gfpga,
		ejection_channels_66__gfpga,
		ejection_channels_65__gfpga,
		ejection_channels_64__gfpga,
		ejection_channels_63__gfpga,
		ejection_channels_62__gfpga,
		ejection_channels_61__gfpga,
		ejection_channels_60__gfpga,
		ejection_channels_59__gfpga,
		ejection_channels_58__gfpga,
		ejection_channels_57__gfpga,
		ejection_channels_56__gfpga,
		ejection_channels_55__gfpga,
		ejection_channels_54__gfpga,
		ejection_channels_53__gfpga,
		ejection_channels_52__gfpga,
		ejection_channels_51__gfpga,
		ejection_channels_50__gfpga,
		ejection_channels_49__gfpga,
		ejection_channels_48__gfpga,
		ejection_channels_47__gfpga,
		ejection_channels_46__gfpga,
		ejection_channels_45__gfpga,
		ejection_channels_44__gfpga,
		ejection_channels_43__gfpga,
		ejection_channels_42__gfpga,
		ejection_channels_41__gfpga,
		ejection_channels_40__gfpga,
		ejection_channels_39__gfpga,
		ejection_channels_38__gfpga,
		ejection_channels_37__gfpga,
		ejection_channels_36__gfpga,
		ejection_channels_35__gfpga,
		ejection_channels_34__gfpga,
		ejection_channels_33__gfpga,
		ejection_channels_32__gfpga,
		ejection_channels_31__gfpga,
		ejection_channels_30__gfpga,
		ejection_channels_29__gfpga,
		ejection_channels_28__gfpga,
		ejection_channels_27__gfpga,
		ejection_channels_26__gfpga,
		ejection_channels_25__gfpga,
		ejection_channels_24__gfpga,
		ejection_channels_23__gfpga,
		ejection_channels_22__gfpga,
		ejection_channels_21__gfpga,
		ejection_channels_20__gfpga,
		ejection_channels_19__gfpga,
		ejection_channels_18__gfpga,
		ejection_channels_17__gfpga,
		ejection_channels_16__gfpga,
		ejection_channels_15__gfpga,
		ejection_channels_14__gfpga,
		ejection_channels_13__gfpga,
		ejection_channels_12__gfpga,
		ejection_channels_11__gfpga,
		ejection_channels_10__gfpga,
		ejection_channels_9__gfpga,
		ejection_channels_8__gfpga,
		ejection_channels_7__gfpga,
		ejection_channels_6__gfpga,
		ejection_channels_5__gfpga,
		ejection_channels_4__gfpga,
		ejection_channels_3__gfpga,
		ejection_channels_2__gfpga,
		ejection_channels_1__gfpga,
		ejection_channels_0__gfpga,
		rtr_error_8__gfpga,
		rtr_error_7__gfpga,
		rtr_error_6__gfpga,
		rtr_error_5__gfpga,
		rtr_error_4__gfpga,
		rtr_error_3__gfpga,
		rtr_error_2__gfpga,
		rtr_error_1__gfpga,
		rtr_error_0__gfpga
	);
// ----- End FPGA Fabric Instanication -------

// ----- Reference Benchmark Instanication -------
	router_mesh REF_DUT(
		clk,
		reset,
		injection_channels_629_,
		injection_channels_628_,
		injection_channels_627_,
		injection_channels_626_,
		injection_channels_625_,
		injection_channels_624_,
		injection_channels_623_,
		injection_channels_622_,
		injection_channels_621_,
		injection_channels_620_,
		injection_channels_619_,
		injection_channels_618_,
		injection_channels_617_,
		injection_channels_616_,
		injection_channels_615_,
		injection_channels_614_,
		injection_channels_613_,
		injection_channels_612_,
		injection_channels_611_,
		injection_channels_610_,
		injection_channels_609_,
		injection_channels_608_,
		injection_channels_607_,
		injection_channels_606_,
		injection_channels_605_,
		injection_channels_604_,
		injection_channels_603_,
		injection_channels_602_,
		injection_channels_601_,
		injection_channels_600_,
		injection_channels_599_,
		injection_channels_598_,
		injection_channels_597_,
		injection_channels_596_,
		injection_channels_595_,
		injection_channels_594_,
		injection_channels_593_,
		injection_channels_592_,
		injection_channels_591_,
		injection_channels_590_,
		injection_channels_589_,
		injection_channels_588_,
		injection_channels_587_,
		injection_channels_586_,
		injection_channels_585_,
		injection_channels_584_,
		injection_channels_583_,
		injection_channels_582_,
		injection_channels_581_,
		injection_channels_580_,
		injection_channels_579_,
		injection_channels_578_,
		injection_channels_577_,
		injection_channels_576_,
		injection_channels_575_,
		injection_channels_574_,
		injection_channels_573_,
		injection_channels_572_,
		injection_channels_571_,
		injection_channels_570_,
		injection_channels_569_,
		injection_channels_568_,
		injection_channels_567_,
		injection_channels_566_,
		injection_channels_565_,
		injection_channels_564_,
		injection_channels_563_,
		injection_channels_562_,
		injection_channels_561_,
		injection_channels_560_,
		injection_channels_559_,
		injection_channels_558_,
		injection_channels_557_,
		injection_channels_556_,
		injection_channels_555_,
		injection_channels_554_,
		injection_channels_553_,
		injection_channels_552_,
		injection_channels_551_,
		injection_channels_550_,
		injection_channels_549_,
		injection_channels_548_,
		injection_channels_547_,
		injection_channels_546_,
		injection_channels_545_,
		injection_channels_544_,
		injection_channels_543_,
		injection_channels_542_,
		injection_channels_541_,
		injection_channels_540_,
		injection_channels_539_,
		injection_channels_538_,
		injection_channels_537_,
		injection_channels_536_,
		injection_channels_535_,
		injection_channels_534_,
		injection_channels_533_,
		injection_channels_532_,
		injection_channels_531_,
		injection_channels_530_,
		injection_channels_529_,
		injection_channels_528_,
		injection_channels_527_,
		injection_channels_526_,
		injection_channels_525_,
		injection_channels_524_,
		injection_channels_523_,
		injection_channels_522_,
		injection_channels_521_,
		injection_channels_520_,
		injection_channels_519_,
		injection_channels_518_,
		injection_channels_517_,
		injection_channels_516_,
		injection_channels_515_,
		injection_channels_514_,
		injection_channels_513_,
		injection_channels_512_,
		injection_channels_511_,
		injection_channels_510_,
		injection_channels_509_,
		injection_channels_508_,
		injection_channels_507_,
		injection_channels_506_,
		injection_channels_505_,
		injection_channels_504_,
		injection_channels_503_,
		injection_channels_502_,
		injection_channels_501_,
		injection_channels_500_,
		injection_channels_499_,
		injection_channels_498_,
		injection_channels_497_,
		injection_channels_496_,
		injection_channels_495_,
		injection_channels_494_,
		injection_channels_493_,
		injection_channels_492_,
		injection_channels_491_,
		injection_channels_490_,
		injection_channels_489_,
		injection_channels_488_,
		injection_channels_487_,
		injection_channels_486_,
		injection_channels_485_,
		injection_channels_484_,
		injection_channels_483_,
		injection_channels_482_,
		injection_channels_481_,
		injection_channels_480_,
		injection_channels_479_,
		injection_channels_478_,
		injection_channels_477_,
		injection_channels_476_,
		injection_channels_475_,
		injection_channels_474_,
		injection_channels_473_,
		injection_channels_472_,
		injection_channels_471_,
		injection_channels_470_,
		injection_channels_469_,
		injection_channels_468_,
		injection_channels_467_,
		injection_channels_466_,
		injection_channels_465_,
		injection_channels_464_,
		injection_channels_463_,
		injection_channels_462_,
		injection_channels_461_,
		injection_channels_460_,
		injection_channels_459_,
		injection_channels_458_,
		injection_channels_457_,
		injection_channels_456_,
		injection_channels_455_,
		injection_channels_454_,
		injection_channels_453_,
		injection_channels_452_,
		injection_channels_451_,
		injection_channels_450_,
		injection_channels_449_,
		injection_channels_448_,
		injection_channels_447_,
		injection_channels_446_,
		injection_channels_445_,
		injection_channels_444_,
		injection_channels_443_,
		injection_channels_442_,
		injection_channels_441_,
		injection_channels_440_,
		injection_channels_439_,
		injection_channels_438_,
		injection_channels_437_,
		injection_channels_436_,
		injection_channels_435_,
		injection_channels_434_,
		injection_channels_433_,
		injection_channels_432_,
		injection_channels_431_,
		injection_channels_430_,
		injection_channels_429_,
		injection_channels_428_,
		injection_channels_427_,
		injection_channels_426_,
		injection_channels_425_,
		injection_channels_424_,
		injection_channels_423_,
		injection_channels_422_,
		injection_channels_421_,
		injection_channels_420_,
		injection_channels_419_,
		injection_channels_418_,
		injection_channels_417_,
		injection_channels_416_,
		injection_channels_415_,
		injection_channels_414_,
		injection_channels_413_,
		injection_channels_412_,
		injection_channels_411_,
		injection_channels_410_,
		injection_channels_409_,
		injection_channels_408_,
		injection_channels_407_,
		injection_channels_406_,
		injection_channels_405_,
		injection_channels_404_,
		injection_channels_403_,
		injection_channels_402_,
		injection_channels_401_,
		injection_channels_400_,
		injection_channels_399_,
		injection_channels_398_,
		injection_channels_397_,
		injection_channels_396_,
		injection_channels_395_,
		injection_channels_394_,
		injection_channels_393_,
		injection_channels_392_,
		injection_channels_391_,
		injection_channels_390_,
		injection_channels_389_,
		injection_channels_388_,
		injection_channels_387_,
		injection_channels_386_,
		injection_channels_385_,
		injection_channels_384_,
		injection_channels_383_,
		injection_channels_382_,
		injection_channels_381_,
		injection_channels_380_,
		injection_channels_379_,
		injection_channels_378_,
		injection_channels_377_,
		injection_channels_376_,
		injection_channels_375_,
		injection_channels_374_,
		injection_channels_373_,
		injection_channels_372_,
		injection_channels_371_,
		injection_channels_370_,
		injection_channels_369_,
		injection_channels_368_,
		injection_channels_367_,
		injection_channels_366_,
		injection_channels_365_,
		injection_channels_364_,
		injection_channels_363_,
		injection_channels_362_,
		injection_channels_361_,
		injection_channels_360_,
		injection_channels_359_,
		injection_channels_358_,
		injection_channels_357_,
		injection_channels_356_,
		injection_channels_355_,
		injection_channels_354_,
		injection_channels_353_,
		injection_channels_352_,
		injection_channels_351_,
		injection_channels_350_,
		injection_channels_349_,
		injection_channels_348_,
		injection_channels_347_,
		injection_channels_346_,
		injection_channels_345_,
		injection_channels_344_,
		injection_channels_343_,
		injection_channels_342_,
		injection_channels_341_,
		injection_channels_340_,
		injection_channels_339_,
		injection_channels_338_,
		injection_channels_337_,
		injection_channels_336_,
		injection_channels_335_,
		injection_channels_334_,
		injection_channels_333_,
		injection_channels_332_,
		injection_channels_331_,
		injection_channels_330_,
		injection_channels_329_,
		injection_channels_328_,
		injection_channels_327_,
		injection_channels_326_,
		injection_channels_325_,
		injection_channels_324_,
		injection_channels_323_,
		injection_channels_322_,
		injection_channels_321_,
		injection_channels_320_,
		injection_channels_319_,
		injection_channels_318_,
		injection_channels_317_,
		injection_channels_316_,
		injection_channels_315_,
		injection_channels_314_,
		injection_channels_313_,
		injection_channels_312_,
		injection_channels_311_,
		injection_channels_310_,
		injection_channels_309_,
		injection_channels_308_,
		injection_channels_307_,
		injection_channels_306_,
		injection_channels_305_,
		injection_channels_304_,
		injection_channels_303_,
		injection_channels_302_,
		injection_channels_301_,
		injection_channels_300_,
		injection_channels_299_,
		injection_channels_298_,
		injection_channels_297_,
		injection_channels_296_,
		injection_channels_295_,
		injection_channels_294_,
		injection_channels_293_,
		injection_channels_292_,
		injection_channels_291_,
		injection_channels_290_,
		injection_channels_289_,
		injection_channels_288_,
		injection_channels_287_,
		injection_channels_286_,
		injection_channels_285_,
		injection_channels_284_,
		injection_channels_283_,
		injection_channels_282_,
		injection_channels_281_,
		injection_channels_280_,
		injection_channels_279_,
		injection_channels_278_,
		injection_channels_277_,
		injection_channels_276_,
		injection_channels_275_,
		injection_channels_274_,
		injection_channels_273_,
		injection_channels_272_,
		injection_channels_271_,
		injection_channels_270_,
		injection_channels_269_,
		injection_channels_268_,
		injection_channels_267_,
		injection_channels_266_,
		injection_channels_265_,
		injection_channels_264_,
		injection_channels_263_,
		injection_channels_262_,
		injection_channels_261_,
		injection_channels_260_,
		injection_channels_259_,
		injection_channels_258_,
		injection_channels_257_,
		injection_channels_256_,
		injection_channels_255_,
		injection_channels_254_,
		injection_channels_253_,
		injection_channels_252_,
		injection_channels_251_,
		injection_channels_250_,
		injection_channels_249_,
		injection_channels_248_,
		injection_channels_247_,
		injection_channels_246_,
		injection_channels_245_,
		injection_channels_244_,
		injection_channels_243_,
		injection_channels_242_,
		injection_channels_241_,
		injection_channels_240_,
		injection_channels_239_,
		injection_channels_238_,
		injection_channels_237_,
		injection_channels_236_,
		injection_channels_235_,
		injection_channels_234_,
		injection_channels_233_,
		injection_channels_232_,
		injection_channels_231_,
		injection_channels_230_,
		injection_channels_229_,
		injection_channels_228_,
		injection_channels_227_,
		injection_channels_226_,
		injection_channels_225_,
		injection_channels_224_,
		injection_channels_223_,
		injection_channels_222_,
		injection_channels_221_,
		injection_channels_220_,
		injection_channels_219_,
		injection_channels_218_,
		injection_channels_217_,
		injection_channels_216_,
		injection_channels_215_,
		injection_channels_214_,
		injection_channels_213_,
		injection_channels_212_,
		injection_channels_211_,
		injection_channels_210_,
		injection_channels_209_,
		injection_channels_208_,
		injection_channels_207_,
		injection_channels_206_,
		injection_channels_205_,
		injection_channels_204_,
		injection_channels_203_,
		injection_channels_202_,
		injection_channels_201_,
		injection_channels_200_,
		injection_channels_199_,
		injection_channels_198_,
		injection_channels_197_,
		injection_channels_196_,
		injection_channels_195_,
		injection_channels_194_,
		injection_channels_193_,
		injection_channels_192_,
		injection_channels_191_,
		injection_channels_190_,
		injection_channels_189_,
		injection_channels_188_,
		injection_channels_187_,
		injection_channels_186_,
		injection_channels_185_,
		injection_channels_184_,
		injection_channels_183_,
		injection_channels_182_,
		injection_channels_181_,
		injection_channels_180_,
		injection_channels_179_,
		injection_channels_178_,
		injection_channels_177_,
		injection_channels_176_,
		injection_channels_175_,
		injection_channels_174_,
		injection_channels_173_,
		injection_channels_172_,
		injection_channels_171_,
		injection_channels_170_,
		injection_channels_169_,
		injection_channels_168_,
		injection_channels_167_,
		injection_channels_166_,
		injection_channels_165_,
		injection_channels_164_,
		injection_channels_163_,
		injection_channels_162_,
		injection_channels_161_,
		injection_channels_160_,
		injection_channels_159_,
		injection_channels_158_,
		injection_channels_157_,
		injection_channels_156_,
		injection_channels_155_,
		injection_channels_154_,
		injection_channels_153_,
		injection_channels_152_,
		injection_channels_151_,
		injection_channels_150_,
		injection_channels_149_,
		injection_channels_148_,
		injection_channels_147_,
		injection_channels_146_,
		injection_channels_145_,
		injection_channels_144_,
		injection_channels_143_,
		injection_channels_142_,
		injection_channels_141_,
		injection_channels_140_,
		injection_channels_139_,
		injection_channels_138_,
		injection_channels_137_,
		injection_channels_136_,
		injection_channels_135_,
		injection_channels_134_,
		injection_channels_133_,
		injection_channels_132_,
		injection_channels_131_,
		injection_channels_130_,
		injection_channels_129_,
		injection_channels_128_,
		injection_channels_127_,
		injection_channels_126_,
		injection_channels_125_,
		injection_channels_124_,
		injection_channels_123_,
		injection_channels_122_,
		injection_channels_121_,
		injection_channels_120_,
		injection_channels_119_,
		injection_channels_118_,
		injection_channels_117_,
		injection_channels_116_,
		injection_channels_115_,
		injection_channels_114_,
		injection_channels_113_,
		injection_channels_112_,
		injection_channels_111_,
		injection_channels_110_,
		injection_channels_109_,
		injection_channels_108_,
		injection_channels_107_,
		injection_channels_106_,
		injection_channels_105_,
		injection_channels_104_,
		injection_channels_103_,
		injection_channels_102_,
		injection_channels_101_,
		injection_channels_100_,
		injection_channels_99_,
		injection_channels_98_,
		injection_channels_97_,
		injection_channels_96_,
		injection_channels_95_,
		injection_channels_94_,
		injection_channels_93_,
		injection_channels_92_,
		injection_channels_91_,
		injection_channels_90_,
		injection_channels_89_,
		injection_channels_88_,
		injection_channels_87_,
		injection_channels_86_,
		injection_channels_85_,
		injection_channels_84_,
		injection_channels_83_,
		injection_channels_82_,
		injection_channels_81_,
		injection_channels_80_,
		injection_channels_79_,
		injection_channels_78_,
		injection_channels_77_,
		injection_channels_76_,
		injection_channels_75_,
		injection_channels_74_,
		injection_channels_73_,
		injection_channels_72_,
		injection_channels_71_,
		injection_channels_70_,
		injection_channels_69_,
		injection_channels_68_,
		injection_channels_67_,
		injection_channels_66_,
		injection_channels_65_,
		injection_channels_64_,
		injection_channels_63_,
		injection_channels_62_,
		injection_channels_61_,
		injection_channels_60_,
		injection_channels_59_,
		injection_channels_58_,
		injection_channels_57_,
		injection_channels_56_,
		injection_channels_55_,
		injection_channels_54_,
		injection_channels_53_,
		injection_channels_52_,
		injection_channels_51_,
		injection_channels_50_,
		injection_channels_49_,
		injection_channels_48_,
		injection_channels_47_,
		injection_channels_46_,
		injection_channels_45_,
		injection_channels_44_,
		injection_channels_43_,
		injection_channels_42_,
		injection_channels_41_,
		injection_channels_40_,
		injection_channels_39_,
		injection_channels_38_,
		injection_channels_37_,
		injection_channels_36_,
		injection_channels_35_,
		injection_channels_34_,
		injection_channels_33_,
		injection_channels_32_,
		injection_channels_31_,
		injection_channels_30_,
		injection_channels_29_,
		injection_channels_28_,
		injection_channels_27_,
		injection_channels_26_,
		injection_channels_25_,
		injection_channels_24_,
		injection_channels_23_,
		injection_channels_22_,
		injection_channels_21_,
		injection_channels_20_,
		injection_channels_19_,
		injection_channels_18_,
		injection_channels_17_,
		injection_channels_16_,
		injection_channels_15_,
		injection_channels_14_,
		injection_channels_13_,
		injection_channels_12_,
		injection_channels_11_,
		injection_channels_10_,
		injection_channels_9_,
		injection_channels_8_,
		injection_channels_7_,
		injection_channels_6_,
		injection_channels_5_,
		injection_channels_4_,
		injection_channels_3_,
		injection_channels_2_,
		injection_channels_1_,
		injection_channels_0_,
		ejection_flow_ctrl_26_,
		ejection_flow_ctrl_25_,
		ejection_flow_ctrl_24_,
		ejection_flow_ctrl_23_,
		ejection_flow_ctrl_22_,
		ejection_flow_ctrl_21_,
		ejection_flow_ctrl_20_,
		ejection_flow_ctrl_19_,
		ejection_flow_ctrl_18_,
		ejection_flow_ctrl_17_,
		ejection_flow_ctrl_16_,
		ejection_flow_ctrl_15_,
		ejection_flow_ctrl_14_,
		ejection_flow_ctrl_13_,
		ejection_flow_ctrl_12_,
		ejection_flow_ctrl_11_,
		ejection_flow_ctrl_10_,
		ejection_flow_ctrl_9_,
		ejection_flow_ctrl_8_,
		ejection_flow_ctrl_7_,
		ejection_flow_ctrl_6_,
		ejection_flow_ctrl_5_,
		ejection_flow_ctrl_4_,
		ejection_flow_ctrl_3_,
		ejection_flow_ctrl_2_,
		ejection_flow_ctrl_1_,
		ejection_flow_ctrl_0_,
		injection_flow_ctrl_26__bench,
		injection_flow_ctrl_25__bench,
		injection_flow_ctrl_24__bench,
		injection_flow_ctrl_23__bench,
		injection_flow_ctrl_22__bench,
		injection_flow_ctrl_21__bench,
		injection_flow_ctrl_20__bench,
		injection_flow_ctrl_19__bench,
		injection_flow_ctrl_18__bench,
		injection_flow_ctrl_17__bench,
		injection_flow_ctrl_16__bench,
		injection_flow_ctrl_15__bench,
		injection_flow_ctrl_14__bench,
		injection_flow_ctrl_13__bench,
		injection_flow_ctrl_12__bench,
		injection_flow_ctrl_11__bench,
		injection_flow_ctrl_10__bench,
		injection_flow_ctrl_9__bench,
		injection_flow_ctrl_8__bench,
		injection_flow_ctrl_7__bench,
		injection_flow_ctrl_6__bench,
		injection_flow_ctrl_5__bench,
		injection_flow_ctrl_4__bench,
		injection_flow_ctrl_3__bench,
		injection_flow_ctrl_2__bench,
		injection_flow_ctrl_1__bench,
		injection_flow_ctrl_0__bench,
		ejection_channels_629__bench,
		ejection_channels_628__bench,
		ejection_channels_627__bench,
		ejection_channels_626__bench,
		ejection_channels_625__bench,
		ejection_channels_624__bench,
		ejection_channels_623__bench,
		ejection_channels_622__bench,
		ejection_channels_621__bench,
		ejection_channels_620__bench,
		ejection_channels_619__bench,
		ejection_channels_618__bench,
		ejection_channels_617__bench,
		ejection_channels_616__bench,
		ejection_channels_615__bench,
		ejection_channels_614__bench,
		ejection_channels_613__bench,
		ejection_channels_612__bench,
		ejection_channels_611__bench,
		ejection_channels_610__bench,
		ejection_channels_609__bench,
		ejection_channels_608__bench,
		ejection_channels_607__bench,
		ejection_channels_606__bench,
		ejection_channels_605__bench,
		ejection_channels_604__bench,
		ejection_channels_603__bench,
		ejection_channels_602__bench,
		ejection_channels_601__bench,
		ejection_channels_600__bench,
		ejection_channels_599__bench,
		ejection_channels_598__bench,
		ejection_channels_597__bench,
		ejection_channels_596__bench,
		ejection_channels_595__bench,
		ejection_channels_594__bench,
		ejection_channels_593__bench,
		ejection_channels_592__bench,
		ejection_channels_591__bench,
		ejection_channels_590__bench,
		ejection_channels_589__bench,
		ejection_channels_588__bench,
		ejection_channels_587__bench,
		ejection_channels_586__bench,
		ejection_channels_585__bench,
		ejection_channels_584__bench,
		ejection_channels_583__bench,
		ejection_channels_582__bench,
		ejection_channels_581__bench,
		ejection_channels_580__bench,
		ejection_channels_579__bench,
		ejection_channels_578__bench,
		ejection_channels_577__bench,
		ejection_channels_576__bench,
		ejection_channels_575__bench,
		ejection_channels_574__bench,
		ejection_channels_573__bench,
		ejection_channels_572__bench,
		ejection_channels_571__bench,
		ejection_channels_570__bench,
		ejection_channels_569__bench,
		ejection_channels_568__bench,
		ejection_channels_567__bench,
		ejection_channels_566__bench,
		ejection_channels_565__bench,
		ejection_channels_564__bench,
		ejection_channels_563__bench,
		ejection_channels_562__bench,
		ejection_channels_561__bench,
		ejection_channels_560__bench,
		ejection_channels_559__bench,
		ejection_channels_558__bench,
		ejection_channels_557__bench,
		ejection_channels_556__bench,
		ejection_channels_555__bench,
		ejection_channels_554__bench,
		ejection_channels_553__bench,
		ejection_channels_552__bench,
		ejection_channels_551__bench,
		ejection_channels_550__bench,
		ejection_channels_549__bench,
		ejection_channels_548__bench,
		ejection_channels_547__bench,
		ejection_channels_546__bench,
		ejection_channels_545__bench,
		ejection_channels_544__bench,
		ejection_channels_543__bench,
		ejection_channels_542__bench,
		ejection_channels_541__bench,
		ejection_channels_540__bench,
		ejection_channels_539__bench,
		ejection_channels_538__bench,
		ejection_channels_537__bench,
		ejection_channels_536__bench,
		ejection_channels_535__bench,
		ejection_channels_534__bench,
		ejection_channels_533__bench,
		ejection_channels_532__bench,
		ejection_channels_531__bench,
		ejection_channels_530__bench,
		ejection_channels_529__bench,
		ejection_channels_528__bench,
		ejection_channels_527__bench,
		ejection_channels_526__bench,
		ejection_channels_525__bench,
		ejection_channels_524__bench,
		ejection_channels_523__bench,
		ejection_channels_522__bench,
		ejection_channels_521__bench,
		ejection_channels_520__bench,
		ejection_channels_519__bench,
		ejection_channels_518__bench,
		ejection_channels_517__bench,
		ejection_channels_516__bench,
		ejection_channels_515__bench,
		ejection_channels_514__bench,
		ejection_channels_513__bench,
		ejection_channels_512__bench,
		ejection_channels_511__bench,
		ejection_channels_510__bench,
		ejection_channels_509__bench,
		ejection_channels_508__bench,
		ejection_channels_507__bench,
		ejection_channels_506__bench,
		ejection_channels_505__bench,
		ejection_channels_504__bench,
		ejection_channels_503__bench,
		ejection_channels_502__bench,
		ejection_channels_501__bench,
		ejection_channels_500__bench,
		ejection_channels_499__bench,
		ejection_channels_498__bench,
		ejection_channels_497__bench,
		ejection_channels_496__bench,
		ejection_channels_495__bench,
		ejection_channels_494__bench,
		ejection_channels_493__bench,
		ejection_channels_492__bench,
		ejection_channels_491__bench,
		ejection_channels_490__bench,
		ejection_channels_489__bench,
		ejection_channels_488__bench,
		ejection_channels_487__bench,
		ejection_channels_486__bench,
		ejection_channels_485__bench,
		ejection_channels_484__bench,
		ejection_channels_483__bench,
		ejection_channels_482__bench,
		ejection_channels_481__bench,
		ejection_channels_480__bench,
		ejection_channels_479__bench,
		ejection_channels_478__bench,
		ejection_channels_477__bench,
		ejection_channels_476__bench,
		ejection_channels_475__bench,
		ejection_channels_474__bench,
		ejection_channels_473__bench,
		ejection_channels_472__bench,
		ejection_channels_471__bench,
		ejection_channels_470__bench,
		ejection_channels_469__bench,
		ejection_channels_468__bench,
		ejection_channels_467__bench,
		ejection_channels_466__bench,
		ejection_channels_465__bench,
		ejection_channels_464__bench,
		ejection_channels_463__bench,
		ejection_channels_462__bench,
		ejection_channels_461__bench,
		ejection_channels_460__bench,
		ejection_channels_459__bench,
		ejection_channels_458__bench,
		ejection_channels_457__bench,
		ejection_channels_456__bench,
		ejection_channels_455__bench,
		ejection_channels_454__bench,
		ejection_channels_453__bench,
		ejection_channels_452__bench,
		ejection_channels_451__bench,
		ejection_channels_450__bench,
		ejection_channels_449__bench,
		ejection_channels_448__bench,
		ejection_channels_447__bench,
		ejection_channels_446__bench,
		ejection_channels_445__bench,
		ejection_channels_444__bench,
		ejection_channels_443__bench,
		ejection_channels_442__bench,
		ejection_channels_441__bench,
		ejection_channels_440__bench,
		ejection_channels_439__bench,
		ejection_channels_438__bench,
		ejection_channels_437__bench,
		ejection_channels_436__bench,
		ejection_channels_435__bench,
		ejection_channels_434__bench,
		ejection_channels_433__bench,
		ejection_channels_432__bench,
		ejection_channels_431__bench,
		ejection_channels_430__bench,
		ejection_channels_429__bench,
		ejection_channels_428__bench,
		ejection_channels_427__bench,
		ejection_channels_426__bench,
		ejection_channels_425__bench,
		ejection_channels_424__bench,
		ejection_channels_423__bench,
		ejection_channels_422__bench,
		ejection_channels_421__bench,
		ejection_channels_420__bench,
		ejection_channels_419__bench,
		ejection_channels_418__bench,
		ejection_channels_417__bench,
		ejection_channels_416__bench,
		ejection_channels_415__bench,
		ejection_channels_414__bench,
		ejection_channels_413__bench,
		ejection_channels_412__bench,
		ejection_channels_411__bench,
		ejection_channels_410__bench,
		ejection_channels_409__bench,
		ejection_channels_408__bench,
		ejection_channels_407__bench,
		ejection_channels_406__bench,
		ejection_channels_405__bench,
		ejection_channels_404__bench,
		ejection_channels_403__bench,
		ejection_channels_402__bench,
		ejection_channels_401__bench,
		ejection_channels_400__bench,
		ejection_channels_399__bench,
		ejection_channels_398__bench,
		ejection_channels_397__bench,
		ejection_channels_396__bench,
		ejection_channels_395__bench,
		ejection_channels_394__bench,
		ejection_channels_393__bench,
		ejection_channels_392__bench,
		ejection_channels_391__bench,
		ejection_channels_390__bench,
		ejection_channels_389__bench,
		ejection_channels_388__bench,
		ejection_channels_387__bench,
		ejection_channels_386__bench,
		ejection_channels_385__bench,
		ejection_channels_384__bench,
		ejection_channels_383__bench,
		ejection_channels_382__bench,
		ejection_channels_381__bench,
		ejection_channels_380__bench,
		ejection_channels_379__bench,
		ejection_channels_378__bench,
		ejection_channels_377__bench,
		ejection_channels_376__bench,
		ejection_channels_375__bench,
		ejection_channels_374__bench,
		ejection_channels_373__bench,
		ejection_channels_372__bench,
		ejection_channels_371__bench,
		ejection_channels_370__bench,
		ejection_channels_369__bench,
		ejection_channels_368__bench,
		ejection_channels_367__bench,
		ejection_channels_366__bench,
		ejection_channels_365__bench,
		ejection_channels_364__bench,
		ejection_channels_363__bench,
		ejection_channels_362__bench,
		ejection_channels_361__bench,
		ejection_channels_360__bench,
		ejection_channels_359__bench,
		ejection_channels_358__bench,
		ejection_channels_357__bench,
		ejection_channels_356__bench,
		ejection_channels_355__bench,
		ejection_channels_354__bench,
		ejection_channels_353__bench,
		ejection_channels_352__bench,
		ejection_channels_351__bench,
		ejection_channels_350__bench,
		ejection_channels_349__bench,
		ejection_channels_348__bench,
		ejection_channels_347__bench,
		ejection_channels_346__bench,
		ejection_channels_345__bench,
		ejection_channels_344__bench,
		ejection_channels_343__bench,
		ejection_channels_342__bench,
		ejection_channels_341__bench,
		ejection_channels_340__bench,
		ejection_channels_339__bench,
		ejection_channels_338__bench,
		ejection_channels_337__bench,
		ejection_channels_336__bench,
		ejection_channels_335__bench,
		ejection_channels_334__bench,
		ejection_channels_333__bench,
		ejection_channels_332__bench,
		ejection_channels_331__bench,
		ejection_channels_330__bench,
		ejection_channels_329__bench,
		ejection_channels_328__bench,
		ejection_channels_327__bench,
		ejection_channels_326__bench,
		ejection_channels_325__bench,
		ejection_channels_324__bench,
		ejection_channels_323__bench,
		ejection_channels_322__bench,
		ejection_channels_321__bench,
		ejection_channels_320__bench,
		ejection_channels_319__bench,
		ejection_channels_318__bench,
		ejection_channels_317__bench,
		ejection_channels_316__bench,
		ejection_channels_315__bench,
		ejection_channels_314__bench,
		ejection_channels_313__bench,
		ejection_channels_312__bench,
		ejection_channels_311__bench,
		ejection_channels_310__bench,
		ejection_channels_309__bench,
		ejection_channels_308__bench,
		ejection_channels_307__bench,
		ejection_channels_306__bench,
		ejection_channels_305__bench,
		ejection_channels_304__bench,
		ejection_channels_303__bench,
		ejection_channels_302__bench,
		ejection_channels_301__bench,
		ejection_channels_300__bench,
		ejection_channels_299__bench,
		ejection_channels_298__bench,
		ejection_channels_297__bench,
		ejection_channels_296__bench,
		ejection_channels_295__bench,
		ejection_channels_294__bench,
		ejection_channels_293__bench,
		ejection_channels_292__bench,
		ejection_channels_291__bench,
		ejection_channels_290__bench,
		ejection_channels_289__bench,
		ejection_channels_288__bench,
		ejection_channels_287__bench,
		ejection_channels_286__bench,
		ejection_channels_285__bench,
		ejection_channels_284__bench,
		ejection_channels_283__bench,
		ejection_channels_282__bench,
		ejection_channels_281__bench,
		ejection_channels_280__bench,
		ejection_channels_279__bench,
		ejection_channels_278__bench,
		ejection_channels_277__bench,
		ejection_channels_276__bench,
		ejection_channels_275__bench,
		ejection_channels_274__bench,
		ejection_channels_273__bench,
		ejection_channels_272__bench,
		ejection_channels_271__bench,
		ejection_channels_270__bench,
		ejection_channels_269__bench,
		ejection_channels_268__bench,
		ejection_channels_267__bench,
		ejection_channels_266__bench,
		ejection_channels_265__bench,
		ejection_channels_264__bench,
		ejection_channels_263__bench,
		ejection_channels_262__bench,
		ejection_channels_261__bench,
		ejection_channels_260__bench,
		ejection_channels_259__bench,
		ejection_channels_258__bench,
		ejection_channels_257__bench,
		ejection_channels_256__bench,
		ejection_channels_255__bench,
		ejection_channels_254__bench,
		ejection_channels_253__bench,
		ejection_channels_252__bench,
		ejection_channels_251__bench,
		ejection_channels_250__bench,
		ejection_channels_249__bench,
		ejection_channels_248__bench,
		ejection_channels_247__bench,
		ejection_channels_246__bench,
		ejection_channels_245__bench,
		ejection_channels_244__bench,
		ejection_channels_243__bench,
		ejection_channels_242__bench,
		ejection_channels_241__bench,
		ejection_channels_240__bench,
		ejection_channels_239__bench,
		ejection_channels_238__bench,
		ejection_channels_237__bench,
		ejection_channels_236__bench,
		ejection_channels_235__bench,
		ejection_channels_234__bench,
		ejection_channels_233__bench,
		ejection_channels_232__bench,
		ejection_channels_231__bench,
		ejection_channels_230__bench,
		ejection_channels_229__bench,
		ejection_channels_228__bench,
		ejection_channels_227__bench,
		ejection_channels_226__bench,
		ejection_channels_225__bench,
		ejection_channels_224__bench,
		ejection_channels_223__bench,
		ejection_channels_222__bench,
		ejection_channels_221__bench,
		ejection_channels_220__bench,
		ejection_channels_219__bench,
		ejection_channels_218__bench,
		ejection_channels_217__bench,
		ejection_channels_216__bench,
		ejection_channels_215__bench,
		ejection_channels_214__bench,
		ejection_channels_213__bench,
		ejection_channels_212__bench,
		ejection_channels_211__bench,
		ejection_channels_210__bench,
		ejection_channels_209__bench,
		ejection_channels_208__bench,
		ejection_channels_207__bench,
		ejection_channels_206__bench,
		ejection_channels_205__bench,
		ejection_channels_204__bench,
		ejection_channels_203__bench,
		ejection_channels_202__bench,
		ejection_channels_201__bench,
		ejection_channels_200__bench,
		ejection_channels_199__bench,
		ejection_channels_198__bench,
		ejection_channels_197__bench,
		ejection_channels_196__bench,
		ejection_channels_195__bench,
		ejection_channels_194__bench,
		ejection_channels_193__bench,
		ejection_channels_192__bench,
		ejection_channels_191__bench,
		ejection_channels_190__bench,
		ejection_channels_189__bench,
		ejection_channels_188__bench,
		ejection_channels_187__bench,
		ejection_channels_186__bench,
		ejection_channels_185__bench,
		ejection_channels_184__bench,
		ejection_channels_183__bench,
		ejection_channels_182__bench,
		ejection_channels_181__bench,
		ejection_channels_180__bench,
		ejection_channels_179__bench,
		ejection_channels_178__bench,
		ejection_channels_177__bench,
		ejection_channels_176__bench,
		ejection_channels_175__bench,
		ejection_channels_174__bench,
		ejection_channels_173__bench,
		ejection_channels_172__bench,
		ejection_channels_171__bench,
		ejection_channels_170__bench,
		ejection_channels_169__bench,
		ejection_channels_168__bench,
		ejection_channels_167__bench,
		ejection_channels_166__bench,
		ejection_channels_165__bench,
		ejection_channels_164__bench,
		ejection_channels_163__bench,
		ejection_channels_162__bench,
		ejection_channels_161__bench,
		ejection_channels_160__bench,
		ejection_channels_159__bench,
		ejection_channels_158__bench,
		ejection_channels_157__bench,
		ejection_channels_156__bench,
		ejection_channels_155__bench,
		ejection_channels_154__bench,
		ejection_channels_153__bench,
		ejection_channels_152__bench,
		ejection_channels_151__bench,
		ejection_channels_150__bench,
		ejection_channels_149__bench,
		ejection_channels_148__bench,
		ejection_channels_147__bench,
		ejection_channels_146__bench,
		ejection_channels_145__bench,
		ejection_channels_144__bench,
		ejection_channels_143__bench,
		ejection_channels_142__bench,
		ejection_channels_141__bench,
		ejection_channels_140__bench,
		ejection_channels_139__bench,
		ejection_channels_138__bench,
		ejection_channels_137__bench,
		ejection_channels_136__bench,
		ejection_channels_135__bench,
		ejection_channels_134__bench,
		ejection_channels_133__bench,
		ejection_channels_132__bench,
		ejection_channels_131__bench,
		ejection_channels_130__bench,
		ejection_channels_129__bench,
		ejection_channels_128__bench,
		ejection_channels_127__bench,
		ejection_channels_126__bench,
		ejection_channels_125__bench,
		ejection_channels_124__bench,
		ejection_channels_123__bench,
		ejection_channels_122__bench,
		ejection_channels_121__bench,
		ejection_channels_120__bench,
		ejection_channels_119__bench,
		ejection_channels_118__bench,
		ejection_channels_117__bench,
		ejection_channels_116__bench,
		ejection_channels_115__bench,
		ejection_channels_114__bench,
		ejection_channels_113__bench,
		ejection_channels_112__bench,
		ejection_channels_111__bench,
		ejection_channels_110__bench,
		ejection_channels_109__bench,
		ejection_channels_108__bench,
		ejection_channels_107__bench,
		ejection_channels_106__bench,
		ejection_channels_105__bench,
		ejection_channels_104__bench,
		ejection_channels_103__bench,
		ejection_channels_102__bench,
		ejection_channels_101__bench,
		ejection_channels_100__bench,
		ejection_channels_99__bench,
		ejection_channels_98__bench,
		ejection_channels_97__bench,
		ejection_channels_96__bench,
		ejection_channels_95__bench,
		ejection_channels_94__bench,
		ejection_channels_93__bench,
		ejection_channels_92__bench,
		ejection_channels_91__bench,
		ejection_channels_90__bench,
		ejection_channels_89__bench,
		ejection_channels_88__bench,
		ejection_channels_87__bench,
		ejection_channels_86__bench,
		ejection_channels_85__bench,
		ejection_channels_84__bench,
		ejection_channels_83__bench,
		ejection_channels_82__bench,
		ejection_channels_81__bench,
		ejection_channels_80__bench,
		ejection_channels_79__bench,
		ejection_channels_78__bench,
		ejection_channels_77__bench,
		ejection_channels_76__bench,
		ejection_channels_75__bench,
		ejection_channels_74__bench,
		ejection_channels_73__bench,
		ejection_channels_72__bench,
		ejection_channels_71__bench,
		ejection_channels_70__bench,
		ejection_channels_69__bench,
		ejection_channels_68__bench,
		ejection_channels_67__bench,
		ejection_channels_66__bench,
		ejection_channels_65__bench,
		ejection_channels_64__bench,
		ejection_channels_63__bench,
		ejection_channels_62__bench,
		ejection_channels_61__bench,
		ejection_channels_60__bench,
		ejection_channels_59__bench,
		ejection_channels_58__bench,
		ejection_channels_57__bench,
		ejection_channels_56__bench,
		ejection_channels_55__bench,
		ejection_channels_54__bench,
		ejection_channels_53__bench,
		ejection_channels_52__bench,
		ejection_channels_51__bench,
		ejection_channels_50__bench,
		ejection_channels_49__bench,
		ejection_channels_48__bench,
		ejection_channels_47__bench,
		ejection_channels_46__bench,
		ejection_channels_45__bench,
		ejection_channels_44__bench,
		ejection_channels_43__bench,
		ejection_channels_42__bench,
		ejection_channels_41__bench,
		ejection_channels_40__bench,
		ejection_channels_39__bench,
		ejection_channels_38__bench,
		ejection_channels_37__bench,
		ejection_channels_36__bench,
		ejection_channels_35__bench,
		ejection_channels_34__bench,
		ejection_channels_33__bench,
		ejection_channels_32__bench,
		ejection_channels_31__bench,
		ejection_channels_30__bench,
		ejection_channels_29__bench,
		ejection_channels_28__bench,
		ejection_channels_27__bench,
		ejection_channels_26__bench,
		ejection_channels_25__bench,
		ejection_channels_24__bench,
		ejection_channels_23__bench,
		ejection_channels_22__bench,
		ejection_channels_21__bench,
		ejection_channels_20__bench,
		ejection_channels_19__bench,
		ejection_channels_18__bench,
		ejection_channels_17__bench,
		ejection_channels_16__bench,
		ejection_channels_15__bench,
		ejection_channels_14__bench,
		ejection_channels_13__bench,
		ejection_channels_12__bench,
		ejection_channels_11__bench,
		ejection_channels_10__bench,
		ejection_channels_9__bench,
		ejection_channels_8__bench,
		ejection_channels_7__bench,
		ejection_channels_6__bench,
		ejection_channels_5__bench,
		ejection_channels_4__bench,
		ejection_channels_3__bench,
		ejection_channels_2__bench,
		ejection_channels_1__bench,
		ejection_channels_0__bench,
		rtr_error_8__bench,
		rtr_error_7__bench,
		rtr_error_6__bench,
		rtr_error_5__bench,
		rtr_error_4__bench,
		rtr_error_3__bench,
		rtr_error_2__bench,
		rtr_error_1__bench,
		rtr_error_0__bench
	);
// ----- End reference Benchmark Instanication -------

// ----- Clock 'clk' Initialization -------
	initial begin
		clk[0] <= 1'b0;
		while(1) begin
			#1
			clk[0] <= !clk[0];
		end
	end

// ----- Begin reset signal generation -----
// ----- End reset signal generation -----

// ----- Input Initialization -------
	initial begin
		reset <= 1'b0;
		injection_channels_629_ <= 1'b0;
		injection_channels_628_ <= 1'b0;
		injection_channels_627_ <= 1'b0;
		injection_channels_626_ <= 1'b0;
		injection_channels_625_ <= 1'b0;
		injection_channels_624_ <= 1'b0;
		injection_channels_623_ <= 1'b0;
		injection_channels_622_ <= 1'b0;
		injection_channels_621_ <= 1'b0;
		injection_channels_620_ <= 1'b0;
		injection_channels_619_ <= 1'b0;
		injection_channels_618_ <= 1'b0;
		injection_channels_617_ <= 1'b0;
		injection_channels_616_ <= 1'b0;
		injection_channels_615_ <= 1'b0;
		injection_channels_614_ <= 1'b0;
		injection_channels_613_ <= 1'b0;
		injection_channels_612_ <= 1'b0;
		injection_channels_611_ <= 1'b0;
		injection_channels_610_ <= 1'b0;
		injection_channels_609_ <= 1'b0;
		injection_channels_608_ <= 1'b0;
		injection_channels_607_ <= 1'b0;
		injection_channels_606_ <= 1'b0;
		injection_channels_605_ <= 1'b0;
		injection_channels_604_ <= 1'b0;
		injection_channels_603_ <= 1'b0;
		injection_channels_602_ <= 1'b0;
		injection_channels_601_ <= 1'b0;
		injection_channels_600_ <= 1'b0;
		injection_channels_599_ <= 1'b0;
		injection_channels_598_ <= 1'b0;
		injection_channels_597_ <= 1'b0;
		injection_channels_596_ <= 1'b0;
		injection_channels_595_ <= 1'b0;
		injection_channels_594_ <= 1'b0;
		injection_channels_593_ <= 1'b0;
		injection_channels_592_ <= 1'b0;
		injection_channels_591_ <= 1'b0;
		injection_channels_590_ <= 1'b0;
		injection_channels_589_ <= 1'b0;
		injection_channels_588_ <= 1'b0;
		injection_channels_587_ <= 1'b0;
		injection_channels_586_ <= 1'b0;
		injection_channels_585_ <= 1'b0;
		injection_channels_584_ <= 1'b0;
		injection_channels_583_ <= 1'b0;
		injection_channels_582_ <= 1'b0;
		injection_channels_581_ <= 1'b0;
		injection_channels_580_ <= 1'b0;
		injection_channels_579_ <= 1'b0;
		injection_channels_578_ <= 1'b0;
		injection_channels_577_ <= 1'b0;
		injection_channels_576_ <= 1'b0;
		injection_channels_575_ <= 1'b0;
		injection_channels_574_ <= 1'b0;
		injection_channels_573_ <= 1'b0;
		injection_channels_572_ <= 1'b0;
		injection_channels_571_ <= 1'b0;
		injection_channels_570_ <= 1'b0;
		injection_channels_569_ <= 1'b0;
		injection_channels_568_ <= 1'b0;
		injection_channels_567_ <= 1'b0;
		injection_channels_566_ <= 1'b0;
		injection_channels_565_ <= 1'b0;
		injection_channels_564_ <= 1'b0;
		injection_channels_563_ <= 1'b0;
		injection_channels_562_ <= 1'b0;
		injection_channels_561_ <= 1'b0;
		injection_channels_560_ <= 1'b0;
		injection_channels_559_ <= 1'b0;
		injection_channels_558_ <= 1'b0;
		injection_channels_557_ <= 1'b0;
		injection_channels_556_ <= 1'b0;
		injection_channels_555_ <= 1'b0;
		injection_channels_554_ <= 1'b0;
		injection_channels_553_ <= 1'b0;
		injection_channels_552_ <= 1'b0;
		injection_channels_551_ <= 1'b0;
		injection_channels_550_ <= 1'b0;
		injection_channels_549_ <= 1'b0;
		injection_channels_548_ <= 1'b0;
		injection_channels_547_ <= 1'b0;
		injection_channels_546_ <= 1'b0;
		injection_channels_545_ <= 1'b0;
		injection_channels_544_ <= 1'b0;
		injection_channels_543_ <= 1'b0;
		injection_channels_542_ <= 1'b0;
		injection_channels_541_ <= 1'b0;
		injection_channels_540_ <= 1'b0;
		injection_channels_539_ <= 1'b0;
		injection_channels_538_ <= 1'b0;
		injection_channels_537_ <= 1'b0;
		injection_channels_536_ <= 1'b0;
		injection_channels_535_ <= 1'b0;
		injection_channels_534_ <= 1'b0;
		injection_channels_533_ <= 1'b0;
		injection_channels_532_ <= 1'b0;
		injection_channels_531_ <= 1'b0;
		injection_channels_530_ <= 1'b0;
		injection_channels_529_ <= 1'b0;
		injection_channels_528_ <= 1'b0;
		injection_channels_527_ <= 1'b0;
		injection_channels_526_ <= 1'b0;
		injection_channels_525_ <= 1'b0;
		injection_channels_524_ <= 1'b0;
		injection_channels_523_ <= 1'b0;
		injection_channels_522_ <= 1'b0;
		injection_channels_521_ <= 1'b0;
		injection_channels_520_ <= 1'b0;
		injection_channels_519_ <= 1'b0;
		injection_channels_518_ <= 1'b0;
		injection_channels_517_ <= 1'b0;
		injection_channels_516_ <= 1'b0;
		injection_channels_515_ <= 1'b0;
		injection_channels_514_ <= 1'b0;
		injection_channels_513_ <= 1'b0;
		injection_channels_512_ <= 1'b0;
		injection_channels_511_ <= 1'b0;
		injection_channels_510_ <= 1'b0;
		injection_channels_509_ <= 1'b0;
		injection_channels_508_ <= 1'b0;
		injection_channels_507_ <= 1'b0;
		injection_channels_506_ <= 1'b0;
		injection_channels_505_ <= 1'b0;
		injection_channels_504_ <= 1'b0;
		injection_channels_503_ <= 1'b0;
		injection_channels_502_ <= 1'b0;
		injection_channels_501_ <= 1'b0;
		injection_channels_500_ <= 1'b0;
		injection_channels_499_ <= 1'b0;
		injection_channels_498_ <= 1'b0;
		injection_channels_497_ <= 1'b0;
		injection_channels_496_ <= 1'b0;
		injection_channels_495_ <= 1'b0;
		injection_channels_494_ <= 1'b0;
		injection_channels_493_ <= 1'b0;
		injection_channels_492_ <= 1'b0;
		injection_channels_491_ <= 1'b0;
		injection_channels_490_ <= 1'b0;
		injection_channels_489_ <= 1'b0;
		injection_channels_488_ <= 1'b0;
		injection_channels_487_ <= 1'b0;
		injection_channels_486_ <= 1'b0;
		injection_channels_485_ <= 1'b0;
		injection_channels_484_ <= 1'b0;
		injection_channels_483_ <= 1'b0;
		injection_channels_482_ <= 1'b0;
		injection_channels_481_ <= 1'b0;
		injection_channels_480_ <= 1'b0;
		injection_channels_479_ <= 1'b0;
		injection_channels_478_ <= 1'b0;
		injection_channels_477_ <= 1'b0;
		injection_channels_476_ <= 1'b0;
		injection_channels_475_ <= 1'b0;
		injection_channels_474_ <= 1'b0;
		injection_channels_473_ <= 1'b0;
		injection_channels_472_ <= 1'b0;
		injection_channels_471_ <= 1'b0;
		injection_channels_470_ <= 1'b0;
		injection_channels_469_ <= 1'b0;
		injection_channels_468_ <= 1'b0;
		injection_channels_467_ <= 1'b0;
		injection_channels_466_ <= 1'b0;
		injection_channels_465_ <= 1'b0;
		injection_channels_464_ <= 1'b0;
		injection_channels_463_ <= 1'b0;
		injection_channels_462_ <= 1'b0;
		injection_channels_461_ <= 1'b0;
		injection_channels_460_ <= 1'b0;
		injection_channels_459_ <= 1'b0;
		injection_channels_458_ <= 1'b0;
		injection_channels_457_ <= 1'b0;
		injection_channels_456_ <= 1'b0;
		injection_channels_455_ <= 1'b0;
		injection_channels_454_ <= 1'b0;
		injection_channels_453_ <= 1'b0;
		injection_channels_452_ <= 1'b0;
		injection_channels_451_ <= 1'b0;
		injection_channels_450_ <= 1'b0;
		injection_channels_449_ <= 1'b0;
		injection_channels_448_ <= 1'b0;
		injection_channels_447_ <= 1'b0;
		injection_channels_446_ <= 1'b0;
		injection_channels_445_ <= 1'b0;
		injection_channels_444_ <= 1'b0;
		injection_channels_443_ <= 1'b0;
		injection_channels_442_ <= 1'b0;
		injection_channels_441_ <= 1'b0;
		injection_channels_440_ <= 1'b0;
		injection_channels_439_ <= 1'b0;
		injection_channels_438_ <= 1'b0;
		injection_channels_437_ <= 1'b0;
		injection_channels_436_ <= 1'b0;
		injection_channels_435_ <= 1'b0;
		injection_channels_434_ <= 1'b0;
		injection_channels_433_ <= 1'b0;
		injection_channels_432_ <= 1'b0;
		injection_channels_431_ <= 1'b0;
		injection_channels_430_ <= 1'b0;
		injection_channels_429_ <= 1'b0;
		injection_channels_428_ <= 1'b0;
		injection_channels_427_ <= 1'b0;
		injection_channels_426_ <= 1'b0;
		injection_channels_425_ <= 1'b0;
		injection_channels_424_ <= 1'b0;
		injection_channels_423_ <= 1'b0;
		injection_channels_422_ <= 1'b0;
		injection_channels_421_ <= 1'b0;
		injection_channels_420_ <= 1'b0;
		injection_channels_419_ <= 1'b0;
		injection_channels_418_ <= 1'b0;
		injection_channels_417_ <= 1'b0;
		injection_channels_416_ <= 1'b0;
		injection_channels_415_ <= 1'b0;
		injection_channels_414_ <= 1'b0;
		injection_channels_413_ <= 1'b0;
		injection_channels_412_ <= 1'b0;
		injection_channels_411_ <= 1'b0;
		injection_channels_410_ <= 1'b0;
		injection_channels_409_ <= 1'b0;
		injection_channels_408_ <= 1'b0;
		injection_channels_407_ <= 1'b0;
		injection_channels_406_ <= 1'b0;
		injection_channels_405_ <= 1'b0;
		injection_channels_404_ <= 1'b0;
		injection_channels_403_ <= 1'b0;
		injection_channels_402_ <= 1'b0;
		injection_channels_401_ <= 1'b0;
		injection_channels_400_ <= 1'b0;
		injection_channels_399_ <= 1'b0;
		injection_channels_398_ <= 1'b0;
		injection_channels_397_ <= 1'b0;
		injection_channels_396_ <= 1'b0;
		injection_channels_395_ <= 1'b0;
		injection_channels_394_ <= 1'b0;
		injection_channels_393_ <= 1'b0;
		injection_channels_392_ <= 1'b0;
		injection_channels_391_ <= 1'b0;
		injection_channels_390_ <= 1'b0;
		injection_channels_389_ <= 1'b0;
		injection_channels_388_ <= 1'b0;
		injection_channels_387_ <= 1'b0;
		injection_channels_386_ <= 1'b0;
		injection_channels_385_ <= 1'b0;
		injection_channels_384_ <= 1'b0;
		injection_channels_383_ <= 1'b0;
		injection_channels_382_ <= 1'b0;
		injection_channels_381_ <= 1'b0;
		injection_channels_380_ <= 1'b0;
		injection_channels_379_ <= 1'b0;
		injection_channels_378_ <= 1'b0;
		injection_channels_377_ <= 1'b0;
		injection_channels_376_ <= 1'b0;
		injection_channels_375_ <= 1'b0;
		injection_channels_374_ <= 1'b0;
		injection_channels_373_ <= 1'b0;
		injection_channels_372_ <= 1'b0;
		injection_channels_371_ <= 1'b0;
		injection_channels_370_ <= 1'b0;
		injection_channels_369_ <= 1'b0;
		injection_channels_368_ <= 1'b0;
		injection_channels_367_ <= 1'b0;
		injection_channels_366_ <= 1'b0;
		injection_channels_365_ <= 1'b0;
		injection_channels_364_ <= 1'b0;
		injection_channels_363_ <= 1'b0;
		injection_channels_362_ <= 1'b0;
		injection_channels_361_ <= 1'b0;
		injection_channels_360_ <= 1'b0;
		injection_channels_359_ <= 1'b0;
		injection_channels_358_ <= 1'b0;
		injection_channels_357_ <= 1'b0;
		injection_channels_356_ <= 1'b0;
		injection_channels_355_ <= 1'b0;
		injection_channels_354_ <= 1'b0;
		injection_channels_353_ <= 1'b0;
		injection_channels_352_ <= 1'b0;
		injection_channels_351_ <= 1'b0;
		injection_channels_350_ <= 1'b0;
		injection_channels_349_ <= 1'b0;
		injection_channels_348_ <= 1'b0;
		injection_channels_347_ <= 1'b0;
		injection_channels_346_ <= 1'b0;
		injection_channels_345_ <= 1'b0;
		injection_channels_344_ <= 1'b0;
		injection_channels_343_ <= 1'b0;
		injection_channels_342_ <= 1'b0;
		injection_channels_341_ <= 1'b0;
		injection_channels_340_ <= 1'b0;
		injection_channels_339_ <= 1'b0;
		injection_channels_338_ <= 1'b0;
		injection_channels_337_ <= 1'b0;
		injection_channels_336_ <= 1'b0;
		injection_channels_335_ <= 1'b0;
		injection_channels_334_ <= 1'b0;
		injection_channels_333_ <= 1'b0;
		injection_channels_332_ <= 1'b0;
		injection_channels_331_ <= 1'b0;
		injection_channels_330_ <= 1'b0;
		injection_channels_329_ <= 1'b0;
		injection_channels_328_ <= 1'b0;
		injection_channels_327_ <= 1'b0;
		injection_channels_326_ <= 1'b0;
		injection_channels_325_ <= 1'b0;
		injection_channels_324_ <= 1'b0;
		injection_channels_323_ <= 1'b0;
		injection_channels_322_ <= 1'b0;
		injection_channels_321_ <= 1'b0;
		injection_channels_320_ <= 1'b0;
		injection_channels_319_ <= 1'b0;
		injection_channels_318_ <= 1'b0;
		injection_channels_317_ <= 1'b0;
		injection_channels_316_ <= 1'b0;
		injection_channels_315_ <= 1'b0;
		injection_channels_314_ <= 1'b0;
		injection_channels_313_ <= 1'b0;
		injection_channels_312_ <= 1'b0;
		injection_channels_311_ <= 1'b0;
		injection_channels_310_ <= 1'b0;
		injection_channels_309_ <= 1'b0;
		injection_channels_308_ <= 1'b0;
		injection_channels_307_ <= 1'b0;
		injection_channels_306_ <= 1'b0;
		injection_channels_305_ <= 1'b0;
		injection_channels_304_ <= 1'b0;
		injection_channels_303_ <= 1'b0;
		injection_channels_302_ <= 1'b0;
		injection_channels_301_ <= 1'b0;
		injection_channels_300_ <= 1'b0;
		injection_channels_299_ <= 1'b0;
		injection_channels_298_ <= 1'b0;
		injection_channels_297_ <= 1'b0;
		injection_channels_296_ <= 1'b0;
		injection_channels_295_ <= 1'b0;
		injection_channels_294_ <= 1'b0;
		injection_channels_293_ <= 1'b0;
		injection_channels_292_ <= 1'b0;
		injection_channels_291_ <= 1'b0;
		injection_channels_290_ <= 1'b0;
		injection_channels_289_ <= 1'b0;
		injection_channels_288_ <= 1'b0;
		injection_channels_287_ <= 1'b0;
		injection_channels_286_ <= 1'b0;
		injection_channels_285_ <= 1'b0;
		injection_channels_284_ <= 1'b0;
		injection_channels_283_ <= 1'b0;
		injection_channels_282_ <= 1'b0;
		injection_channels_281_ <= 1'b0;
		injection_channels_280_ <= 1'b0;
		injection_channels_279_ <= 1'b0;
		injection_channels_278_ <= 1'b0;
		injection_channels_277_ <= 1'b0;
		injection_channels_276_ <= 1'b0;
		injection_channels_275_ <= 1'b0;
		injection_channels_274_ <= 1'b0;
		injection_channels_273_ <= 1'b0;
		injection_channels_272_ <= 1'b0;
		injection_channels_271_ <= 1'b0;
		injection_channels_270_ <= 1'b0;
		injection_channels_269_ <= 1'b0;
		injection_channels_268_ <= 1'b0;
		injection_channels_267_ <= 1'b0;
		injection_channels_266_ <= 1'b0;
		injection_channels_265_ <= 1'b0;
		injection_channels_264_ <= 1'b0;
		injection_channels_263_ <= 1'b0;
		injection_channels_262_ <= 1'b0;
		injection_channels_261_ <= 1'b0;
		injection_channels_260_ <= 1'b0;
		injection_channels_259_ <= 1'b0;
		injection_channels_258_ <= 1'b0;
		injection_channels_257_ <= 1'b0;
		injection_channels_256_ <= 1'b0;
		injection_channels_255_ <= 1'b0;
		injection_channels_254_ <= 1'b0;
		injection_channels_253_ <= 1'b0;
		injection_channels_252_ <= 1'b0;
		injection_channels_251_ <= 1'b0;
		injection_channels_250_ <= 1'b0;
		injection_channels_249_ <= 1'b0;
		injection_channels_248_ <= 1'b0;
		injection_channels_247_ <= 1'b0;
		injection_channels_246_ <= 1'b0;
		injection_channels_245_ <= 1'b0;
		injection_channels_244_ <= 1'b0;
		injection_channels_243_ <= 1'b0;
		injection_channels_242_ <= 1'b0;
		injection_channels_241_ <= 1'b0;
		injection_channels_240_ <= 1'b0;
		injection_channels_239_ <= 1'b0;
		injection_channels_238_ <= 1'b0;
		injection_channels_237_ <= 1'b0;
		injection_channels_236_ <= 1'b0;
		injection_channels_235_ <= 1'b0;
		injection_channels_234_ <= 1'b0;
		injection_channels_233_ <= 1'b0;
		injection_channels_232_ <= 1'b0;
		injection_channels_231_ <= 1'b0;
		injection_channels_230_ <= 1'b0;
		injection_channels_229_ <= 1'b0;
		injection_channels_228_ <= 1'b0;
		injection_channels_227_ <= 1'b0;
		injection_channels_226_ <= 1'b0;
		injection_channels_225_ <= 1'b0;
		injection_channels_224_ <= 1'b0;
		injection_channels_223_ <= 1'b0;
		injection_channels_222_ <= 1'b0;
		injection_channels_221_ <= 1'b0;
		injection_channels_220_ <= 1'b0;
		injection_channels_219_ <= 1'b0;
		injection_channels_218_ <= 1'b0;
		injection_channels_217_ <= 1'b0;
		injection_channels_216_ <= 1'b0;
		injection_channels_215_ <= 1'b0;
		injection_channels_214_ <= 1'b0;
		injection_channels_213_ <= 1'b0;
		injection_channels_212_ <= 1'b0;
		injection_channels_211_ <= 1'b0;
		injection_channels_210_ <= 1'b0;
		injection_channels_209_ <= 1'b0;
		injection_channels_208_ <= 1'b0;
		injection_channels_207_ <= 1'b0;
		injection_channels_206_ <= 1'b0;
		injection_channels_205_ <= 1'b0;
		injection_channels_204_ <= 1'b0;
		injection_channels_203_ <= 1'b0;
		injection_channels_202_ <= 1'b0;
		injection_channels_201_ <= 1'b0;
		injection_channels_200_ <= 1'b0;
		injection_channels_199_ <= 1'b0;
		injection_channels_198_ <= 1'b0;
		injection_channels_197_ <= 1'b0;
		injection_channels_196_ <= 1'b0;
		injection_channels_195_ <= 1'b0;
		injection_channels_194_ <= 1'b0;
		injection_channels_193_ <= 1'b0;
		injection_channels_192_ <= 1'b0;
		injection_channels_191_ <= 1'b0;
		injection_channels_190_ <= 1'b0;
		injection_channels_189_ <= 1'b0;
		injection_channels_188_ <= 1'b0;
		injection_channels_187_ <= 1'b0;
		injection_channels_186_ <= 1'b0;
		injection_channels_185_ <= 1'b0;
		injection_channels_184_ <= 1'b0;
		injection_channels_183_ <= 1'b0;
		injection_channels_182_ <= 1'b0;
		injection_channels_181_ <= 1'b0;
		injection_channels_180_ <= 1'b0;
		injection_channels_179_ <= 1'b0;
		injection_channels_178_ <= 1'b0;
		injection_channels_177_ <= 1'b0;
		injection_channels_176_ <= 1'b0;
		injection_channels_175_ <= 1'b0;
		injection_channels_174_ <= 1'b0;
		injection_channels_173_ <= 1'b0;
		injection_channels_172_ <= 1'b0;
		injection_channels_171_ <= 1'b0;
		injection_channels_170_ <= 1'b0;
		injection_channels_169_ <= 1'b0;
		injection_channels_168_ <= 1'b0;
		injection_channels_167_ <= 1'b0;
		injection_channels_166_ <= 1'b0;
		injection_channels_165_ <= 1'b0;
		injection_channels_164_ <= 1'b0;
		injection_channels_163_ <= 1'b0;
		injection_channels_162_ <= 1'b0;
		injection_channels_161_ <= 1'b0;
		injection_channels_160_ <= 1'b0;
		injection_channels_159_ <= 1'b0;
		injection_channels_158_ <= 1'b0;
		injection_channels_157_ <= 1'b0;
		injection_channels_156_ <= 1'b0;
		injection_channels_155_ <= 1'b0;
		injection_channels_154_ <= 1'b0;
		injection_channels_153_ <= 1'b0;
		injection_channels_152_ <= 1'b0;
		injection_channels_151_ <= 1'b0;
		injection_channels_150_ <= 1'b0;
		injection_channels_149_ <= 1'b0;
		injection_channels_148_ <= 1'b0;
		injection_channels_147_ <= 1'b0;
		injection_channels_146_ <= 1'b0;
		injection_channels_145_ <= 1'b0;
		injection_channels_144_ <= 1'b0;
		injection_channels_143_ <= 1'b0;
		injection_channels_142_ <= 1'b0;
		injection_channels_141_ <= 1'b0;
		injection_channels_140_ <= 1'b0;
		injection_channels_139_ <= 1'b0;
		injection_channels_138_ <= 1'b0;
		injection_channels_137_ <= 1'b0;
		injection_channels_136_ <= 1'b0;
		injection_channels_135_ <= 1'b0;
		injection_channels_134_ <= 1'b0;
		injection_channels_133_ <= 1'b0;
		injection_channels_132_ <= 1'b0;
		injection_channels_131_ <= 1'b0;
		injection_channels_130_ <= 1'b0;
		injection_channels_129_ <= 1'b0;
		injection_channels_128_ <= 1'b0;
		injection_channels_127_ <= 1'b0;
		injection_channels_126_ <= 1'b0;
		injection_channels_125_ <= 1'b0;
		injection_channels_124_ <= 1'b0;
		injection_channels_123_ <= 1'b0;
		injection_channels_122_ <= 1'b0;
		injection_channels_121_ <= 1'b0;
		injection_channels_120_ <= 1'b0;
		injection_channels_119_ <= 1'b0;
		injection_channels_118_ <= 1'b0;
		injection_channels_117_ <= 1'b0;
		injection_channels_116_ <= 1'b0;
		injection_channels_115_ <= 1'b0;
		injection_channels_114_ <= 1'b0;
		injection_channels_113_ <= 1'b0;
		injection_channels_112_ <= 1'b0;
		injection_channels_111_ <= 1'b0;
		injection_channels_110_ <= 1'b0;
		injection_channels_109_ <= 1'b0;
		injection_channels_108_ <= 1'b0;
		injection_channels_107_ <= 1'b0;
		injection_channels_106_ <= 1'b0;
		injection_channels_105_ <= 1'b0;
		injection_channels_104_ <= 1'b0;
		injection_channels_103_ <= 1'b0;
		injection_channels_102_ <= 1'b0;
		injection_channels_101_ <= 1'b0;
		injection_channels_100_ <= 1'b0;
		injection_channels_99_ <= 1'b0;
		injection_channels_98_ <= 1'b0;
		injection_channels_97_ <= 1'b0;
		injection_channels_96_ <= 1'b0;
		injection_channels_95_ <= 1'b0;
		injection_channels_94_ <= 1'b0;
		injection_channels_93_ <= 1'b0;
		injection_channels_92_ <= 1'b0;
		injection_channels_91_ <= 1'b0;
		injection_channels_90_ <= 1'b0;
		injection_channels_89_ <= 1'b0;
		injection_channels_88_ <= 1'b0;
		injection_channels_87_ <= 1'b0;
		injection_channels_86_ <= 1'b0;
		injection_channels_85_ <= 1'b0;
		injection_channels_84_ <= 1'b0;
		injection_channels_83_ <= 1'b0;
		injection_channels_82_ <= 1'b0;
		injection_channels_81_ <= 1'b0;
		injection_channels_80_ <= 1'b0;
		injection_channels_79_ <= 1'b0;
		injection_channels_78_ <= 1'b0;
		injection_channels_77_ <= 1'b0;
		injection_channels_76_ <= 1'b0;
		injection_channels_75_ <= 1'b0;
		injection_channels_74_ <= 1'b0;
		injection_channels_73_ <= 1'b0;
		injection_channels_72_ <= 1'b0;
		injection_channels_71_ <= 1'b0;
		injection_channels_70_ <= 1'b0;
		injection_channels_69_ <= 1'b0;
		injection_channels_68_ <= 1'b0;
		injection_channels_67_ <= 1'b0;
		injection_channels_66_ <= 1'b0;
		injection_channels_65_ <= 1'b0;
		injection_channels_64_ <= 1'b0;
		injection_channels_63_ <= 1'b0;
		injection_channels_62_ <= 1'b0;
		injection_channels_61_ <= 1'b0;
		injection_channels_60_ <= 1'b0;
		injection_channels_59_ <= 1'b0;
		injection_channels_58_ <= 1'b0;
		injection_channels_57_ <= 1'b0;
		injection_channels_56_ <= 1'b0;
		injection_channels_55_ <= 1'b0;
		injection_channels_54_ <= 1'b0;
		injection_channels_53_ <= 1'b0;
		injection_channels_52_ <= 1'b0;
		injection_channels_51_ <= 1'b0;
		injection_channels_50_ <= 1'b0;
		injection_channels_49_ <= 1'b0;
		injection_channels_48_ <= 1'b0;
		injection_channels_47_ <= 1'b0;
		injection_channels_46_ <= 1'b0;
		injection_channels_45_ <= 1'b0;
		injection_channels_44_ <= 1'b0;
		injection_channels_43_ <= 1'b0;
		injection_channels_42_ <= 1'b0;
		injection_channels_41_ <= 1'b0;
		injection_channels_40_ <= 1'b0;
		injection_channels_39_ <= 1'b0;
		injection_channels_38_ <= 1'b0;
		injection_channels_37_ <= 1'b0;
		injection_channels_36_ <= 1'b0;
		injection_channels_35_ <= 1'b0;
		injection_channels_34_ <= 1'b0;
		injection_channels_33_ <= 1'b0;
		injection_channels_32_ <= 1'b0;
		injection_channels_31_ <= 1'b0;
		injection_channels_30_ <= 1'b0;
		injection_channels_29_ <= 1'b0;
		injection_channels_28_ <= 1'b0;
		injection_channels_27_ <= 1'b0;
		injection_channels_26_ <= 1'b0;
		injection_channels_25_ <= 1'b0;
		injection_channels_24_ <= 1'b0;
		injection_channels_23_ <= 1'b0;
		injection_channels_22_ <= 1'b0;
		injection_channels_21_ <= 1'b0;
		injection_channels_20_ <= 1'b0;
		injection_channels_19_ <= 1'b0;
		injection_channels_18_ <= 1'b0;
		injection_channels_17_ <= 1'b0;
		injection_channels_16_ <= 1'b0;
		injection_channels_15_ <= 1'b0;
		injection_channels_14_ <= 1'b0;
		injection_channels_13_ <= 1'b0;
		injection_channels_12_ <= 1'b0;
		injection_channels_11_ <= 1'b0;
		injection_channels_10_ <= 1'b0;
		injection_channels_9_ <= 1'b0;
		injection_channels_8_ <= 1'b0;
		injection_channels_7_ <= 1'b0;
		injection_channels_6_ <= 1'b0;
		injection_channels_5_ <= 1'b0;
		injection_channels_4_ <= 1'b0;
		injection_channels_3_ <= 1'b0;
		injection_channels_2_ <= 1'b0;
		injection_channels_1_ <= 1'b0;
		injection_channels_0_ <= 1'b0;
		ejection_flow_ctrl_26_ <= 1'b0;
		ejection_flow_ctrl_25_ <= 1'b0;
		ejection_flow_ctrl_24_ <= 1'b0;
		ejection_flow_ctrl_23_ <= 1'b0;
		ejection_flow_ctrl_22_ <= 1'b0;
		ejection_flow_ctrl_21_ <= 1'b0;
		ejection_flow_ctrl_20_ <= 1'b0;
		ejection_flow_ctrl_19_ <= 1'b0;
		ejection_flow_ctrl_18_ <= 1'b0;
		ejection_flow_ctrl_17_ <= 1'b0;
		ejection_flow_ctrl_16_ <= 1'b0;
		ejection_flow_ctrl_15_ <= 1'b0;
		ejection_flow_ctrl_14_ <= 1'b0;
		ejection_flow_ctrl_13_ <= 1'b0;
		ejection_flow_ctrl_12_ <= 1'b0;
		ejection_flow_ctrl_11_ <= 1'b0;
		ejection_flow_ctrl_10_ <= 1'b0;
		ejection_flow_ctrl_9_ <= 1'b0;
		ejection_flow_ctrl_8_ <= 1'b0;
		ejection_flow_ctrl_7_ <= 1'b0;
		ejection_flow_ctrl_6_ <= 1'b0;
		ejection_flow_ctrl_5_ <= 1'b0;
		ejection_flow_ctrl_4_ <= 1'b0;
		ejection_flow_ctrl_3_ <= 1'b0;
		ejection_flow_ctrl_2_ <= 1'b0;
		ejection_flow_ctrl_1_ <= 1'b0;
		ejection_flow_ctrl_0_ <= 1'b0;

		injection_flow_ctrl_26__flag[0] <= 1'b0;
		injection_flow_ctrl_25__flag[0] <= 1'b0;
		injection_flow_ctrl_24__flag[0] <= 1'b0;
		injection_flow_ctrl_23__flag[0] <= 1'b0;
		injection_flow_ctrl_22__flag[0] <= 1'b0;
		injection_flow_ctrl_21__flag[0] <= 1'b0;
		injection_flow_ctrl_20__flag[0] <= 1'b0;
		injection_flow_ctrl_19__flag[0] <= 1'b0;
		injection_flow_ctrl_18__flag[0] <= 1'b0;
		injection_flow_ctrl_17__flag[0] <= 1'b0;
		injection_flow_ctrl_16__flag[0] <= 1'b0;
		injection_flow_ctrl_15__flag[0] <= 1'b0;
		injection_flow_ctrl_14__flag[0] <= 1'b0;
		injection_flow_ctrl_13__flag[0] <= 1'b0;
		injection_flow_ctrl_12__flag[0] <= 1'b0;
		injection_flow_ctrl_11__flag[0] <= 1'b0;
		injection_flow_ctrl_10__flag[0] <= 1'b0;
		injection_flow_ctrl_9__flag[0] <= 1'b0;
		injection_flow_ctrl_8__flag[0] <= 1'b0;
		injection_flow_ctrl_7__flag[0] <= 1'b0;
		injection_flow_ctrl_6__flag[0] <= 1'b0;
		injection_flow_ctrl_5__flag[0] <= 1'b0;
		injection_flow_ctrl_4__flag[0] <= 1'b0;
		injection_flow_ctrl_3__flag[0] <= 1'b0;
		injection_flow_ctrl_2__flag[0] <= 1'b0;
		injection_flow_ctrl_1__flag[0] <= 1'b0;
		injection_flow_ctrl_0__flag[0] <= 1'b0;
		ejection_channels_629__flag[0] <= 1'b0;
		ejection_channels_628__flag[0] <= 1'b0;
		ejection_channels_627__flag[0] <= 1'b0;
		ejection_channels_626__flag[0] <= 1'b0;
		ejection_channels_625__flag[0] <= 1'b0;
		ejection_channels_624__flag[0] <= 1'b0;
		ejection_channels_623__flag[0] <= 1'b0;
		ejection_channels_622__flag[0] <= 1'b0;
		ejection_channels_621__flag[0] <= 1'b0;
		ejection_channels_620__flag[0] <= 1'b0;
		ejection_channels_619__flag[0] <= 1'b0;
		ejection_channels_618__flag[0] <= 1'b0;
		ejection_channels_617__flag[0] <= 1'b0;
		ejection_channels_616__flag[0] <= 1'b0;
		ejection_channels_615__flag[0] <= 1'b0;
		ejection_channels_614__flag[0] <= 1'b0;
		ejection_channels_613__flag[0] <= 1'b0;
		ejection_channels_612__flag[0] <= 1'b0;
		ejection_channels_611__flag[0] <= 1'b0;
		ejection_channels_610__flag[0] <= 1'b0;
		ejection_channels_609__flag[0] <= 1'b0;
		ejection_channels_608__flag[0] <= 1'b0;
		ejection_channels_607__flag[0] <= 1'b0;
		ejection_channels_606__flag[0] <= 1'b0;
		ejection_channels_605__flag[0] <= 1'b0;
		ejection_channels_604__flag[0] <= 1'b0;
		ejection_channels_603__flag[0] <= 1'b0;
		ejection_channels_602__flag[0] <= 1'b0;
		ejection_channels_601__flag[0] <= 1'b0;
		ejection_channels_600__flag[0] <= 1'b0;
		ejection_channels_599__flag[0] <= 1'b0;
		ejection_channels_598__flag[0] <= 1'b0;
		ejection_channels_597__flag[0] <= 1'b0;
		ejection_channels_596__flag[0] <= 1'b0;
		ejection_channels_595__flag[0] <= 1'b0;
		ejection_channels_594__flag[0] <= 1'b0;
		ejection_channels_593__flag[0] <= 1'b0;
		ejection_channels_592__flag[0] <= 1'b0;
		ejection_channels_591__flag[0] <= 1'b0;
		ejection_channels_590__flag[0] <= 1'b0;
		ejection_channels_589__flag[0] <= 1'b0;
		ejection_channels_588__flag[0] <= 1'b0;
		ejection_channels_587__flag[0] <= 1'b0;
		ejection_channels_586__flag[0] <= 1'b0;
		ejection_channels_585__flag[0] <= 1'b0;
		ejection_channels_584__flag[0] <= 1'b0;
		ejection_channels_583__flag[0] <= 1'b0;
		ejection_channels_582__flag[0] <= 1'b0;
		ejection_channels_581__flag[0] <= 1'b0;
		ejection_channels_580__flag[0] <= 1'b0;
		ejection_channels_579__flag[0] <= 1'b0;
		ejection_channels_578__flag[0] <= 1'b0;
		ejection_channels_577__flag[0] <= 1'b0;
		ejection_channels_576__flag[0] <= 1'b0;
		ejection_channels_575__flag[0] <= 1'b0;
		ejection_channels_574__flag[0] <= 1'b0;
		ejection_channels_573__flag[0] <= 1'b0;
		ejection_channels_572__flag[0] <= 1'b0;
		ejection_channels_571__flag[0] <= 1'b0;
		ejection_channels_570__flag[0] <= 1'b0;
		ejection_channels_569__flag[0] <= 1'b0;
		ejection_channels_568__flag[0] <= 1'b0;
		ejection_channels_567__flag[0] <= 1'b0;
		ejection_channels_566__flag[0] <= 1'b0;
		ejection_channels_565__flag[0] <= 1'b0;
		ejection_channels_564__flag[0] <= 1'b0;
		ejection_channels_563__flag[0] <= 1'b0;
		ejection_channels_562__flag[0] <= 1'b0;
		ejection_channels_561__flag[0] <= 1'b0;
		ejection_channels_560__flag[0] <= 1'b0;
		ejection_channels_559__flag[0] <= 1'b0;
		ejection_channels_558__flag[0] <= 1'b0;
		ejection_channels_557__flag[0] <= 1'b0;
		ejection_channels_556__flag[0] <= 1'b0;
		ejection_channels_555__flag[0] <= 1'b0;
		ejection_channels_554__flag[0] <= 1'b0;
		ejection_channels_553__flag[0] <= 1'b0;
		ejection_channels_552__flag[0] <= 1'b0;
		ejection_channels_551__flag[0] <= 1'b0;
		ejection_channels_550__flag[0] <= 1'b0;
		ejection_channels_549__flag[0] <= 1'b0;
		ejection_channels_548__flag[0] <= 1'b0;
		ejection_channels_547__flag[0] <= 1'b0;
		ejection_channels_546__flag[0] <= 1'b0;
		ejection_channels_545__flag[0] <= 1'b0;
		ejection_channels_544__flag[0] <= 1'b0;
		ejection_channels_543__flag[0] <= 1'b0;
		ejection_channels_542__flag[0] <= 1'b0;
		ejection_channels_541__flag[0] <= 1'b0;
		ejection_channels_540__flag[0] <= 1'b0;
		ejection_channels_539__flag[0] <= 1'b0;
		ejection_channels_538__flag[0] <= 1'b0;
		ejection_channels_537__flag[0] <= 1'b0;
		ejection_channels_536__flag[0] <= 1'b0;
		ejection_channels_535__flag[0] <= 1'b0;
		ejection_channels_534__flag[0] <= 1'b0;
		ejection_channels_533__flag[0] <= 1'b0;
		ejection_channels_532__flag[0] <= 1'b0;
		ejection_channels_531__flag[0] <= 1'b0;
		ejection_channels_530__flag[0] <= 1'b0;
		ejection_channels_529__flag[0] <= 1'b0;
		ejection_channels_528__flag[0] <= 1'b0;
		ejection_channels_527__flag[0] <= 1'b0;
		ejection_channels_526__flag[0] <= 1'b0;
		ejection_channels_525__flag[0] <= 1'b0;
		ejection_channels_524__flag[0] <= 1'b0;
		ejection_channels_523__flag[0] <= 1'b0;
		ejection_channels_522__flag[0] <= 1'b0;
		ejection_channels_521__flag[0] <= 1'b0;
		ejection_channels_520__flag[0] <= 1'b0;
		ejection_channels_519__flag[0] <= 1'b0;
		ejection_channels_518__flag[0] <= 1'b0;
		ejection_channels_517__flag[0] <= 1'b0;
		ejection_channels_516__flag[0] <= 1'b0;
		ejection_channels_515__flag[0] <= 1'b0;
		ejection_channels_514__flag[0] <= 1'b0;
		ejection_channels_513__flag[0] <= 1'b0;
		ejection_channels_512__flag[0] <= 1'b0;
		ejection_channels_511__flag[0] <= 1'b0;
		ejection_channels_510__flag[0] <= 1'b0;
		ejection_channels_509__flag[0] <= 1'b0;
		ejection_channels_508__flag[0] <= 1'b0;
		ejection_channels_507__flag[0] <= 1'b0;
		ejection_channels_506__flag[0] <= 1'b0;
		ejection_channels_505__flag[0] <= 1'b0;
		ejection_channels_504__flag[0] <= 1'b0;
		ejection_channels_503__flag[0] <= 1'b0;
		ejection_channels_502__flag[0] <= 1'b0;
		ejection_channels_501__flag[0] <= 1'b0;
		ejection_channels_500__flag[0] <= 1'b0;
		ejection_channels_499__flag[0] <= 1'b0;
		ejection_channels_498__flag[0] <= 1'b0;
		ejection_channels_497__flag[0] <= 1'b0;
		ejection_channels_496__flag[0] <= 1'b0;
		ejection_channels_495__flag[0] <= 1'b0;
		ejection_channels_494__flag[0] <= 1'b0;
		ejection_channels_493__flag[0] <= 1'b0;
		ejection_channels_492__flag[0] <= 1'b0;
		ejection_channels_491__flag[0] <= 1'b0;
		ejection_channels_490__flag[0] <= 1'b0;
		ejection_channels_489__flag[0] <= 1'b0;
		ejection_channels_488__flag[0] <= 1'b0;
		ejection_channels_487__flag[0] <= 1'b0;
		ejection_channels_486__flag[0] <= 1'b0;
		ejection_channels_485__flag[0] <= 1'b0;
		ejection_channels_484__flag[0] <= 1'b0;
		ejection_channels_483__flag[0] <= 1'b0;
		ejection_channels_482__flag[0] <= 1'b0;
		ejection_channels_481__flag[0] <= 1'b0;
		ejection_channels_480__flag[0] <= 1'b0;
		ejection_channels_479__flag[0] <= 1'b0;
		ejection_channels_478__flag[0] <= 1'b0;
		ejection_channels_477__flag[0] <= 1'b0;
		ejection_channels_476__flag[0] <= 1'b0;
		ejection_channels_475__flag[0] <= 1'b0;
		ejection_channels_474__flag[0] <= 1'b0;
		ejection_channels_473__flag[0] <= 1'b0;
		ejection_channels_472__flag[0] <= 1'b0;
		ejection_channels_471__flag[0] <= 1'b0;
		ejection_channels_470__flag[0] <= 1'b0;
		ejection_channels_469__flag[0] <= 1'b0;
		ejection_channels_468__flag[0] <= 1'b0;
		ejection_channels_467__flag[0] <= 1'b0;
		ejection_channels_466__flag[0] <= 1'b0;
		ejection_channels_465__flag[0] <= 1'b0;
		ejection_channels_464__flag[0] <= 1'b0;
		ejection_channels_463__flag[0] <= 1'b0;
		ejection_channels_462__flag[0] <= 1'b0;
		ejection_channels_461__flag[0] <= 1'b0;
		ejection_channels_460__flag[0] <= 1'b0;
		ejection_channels_459__flag[0] <= 1'b0;
		ejection_channels_458__flag[0] <= 1'b0;
		ejection_channels_457__flag[0] <= 1'b0;
		ejection_channels_456__flag[0] <= 1'b0;
		ejection_channels_455__flag[0] <= 1'b0;
		ejection_channels_454__flag[0] <= 1'b0;
		ejection_channels_453__flag[0] <= 1'b0;
		ejection_channels_452__flag[0] <= 1'b0;
		ejection_channels_451__flag[0] <= 1'b0;
		ejection_channels_450__flag[0] <= 1'b0;
		ejection_channels_449__flag[0] <= 1'b0;
		ejection_channels_448__flag[0] <= 1'b0;
		ejection_channels_447__flag[0] <= 1'b0;
		ejection_channels_446__flag[0] <= 1'b0;
		ejection_channels_445__flag[0] <= 1'b0;
		ejection_channels_444__flag[0] <= 1'b0;
		ejection_channels_443__flag[0] <= 1'b0;
		ejection_channels_442__flag[0] <= 1'b0;
		ejection_channels_441__flag[0] <= 1'b0;
		ejection_channels_440__flag[0] <= 1'b0;
		ejection_channels_439__flag[0] <= 1'b0;
		ejection_channels_438__flag[0] <= 1'b0;
		ejection_channels_437__flag[0] <= 1'b0;
		ejection_channels_436__flag[0] <= 1'b0;
		ejection_channels_435__flag[0] <= 1'b0;
		ejection_channels_434__flag[0] <= 1'b0;
		ejection_channels_433__flag[0] <= 1'b0;
		ejection_channels_432__flag[0] <= 1'b0;
		ejection_channels_431__flag[0] <= 1'b0;
		ejection_channels_430__flag[0] <= 1'b0;
		ejection_channels_429__flag[0] <= 1'b0;
		ejection_channels_428__flag[0] <= 1'b0;
		ejection_channels_427__flag[0] <= 1'b0;
		ejection_channels_426__flag[0] <= 1'b0;
		ejection_channels_425__flag[0] <= 1'b0;
		ejection_channels_424__flag[0] <= 1'b0;
		ejection_channels_423__flag[0] <= 1'b0;
		ejection_channels_422__flag[0] <= 1'b0;
		ejection_channels_421__flag[0] <= 1'b0;
		ejection_channels_420__flag[0] <= 1'b0;
		ejection_channels_419__flag[0] <= 1'b0;
		ejection_channels_418__flag[0] <= 1'b0;
		ejection_channels_417__flag[0] <= 1'b0;
		ejection_channels_416__flag[0] <= 1'b0;
		ejection_channels_415__flag[0] <= 1'b0;
		ejection_channels_414__flag[0] <= 1'b0;
		ejection_channels_413__flag[0] <= 1'b0;
		ejection_channels_412__flag[0] <= 1'b0;
		ejection_channels_411__flag[0] <= 1'b0;
		ejection_channels_410__flag[0] <= 1'b0;
		ejection_channels_409__flag[0] <= 1'b0;
		ejection_channels_408__flag[0] <= 1'b0;
		ejection_channels_407__flag[0] <= 1'b0;
		ejection_channels_406__flag[0] <= 1'b0;
		ejection_channels_405__flag[0] <= 1'b0;
		ejection_channels_404__flag[0] <= 1'b0;
		ejection_channels_403__flag[0] <= 1'b0;
		ejection_channels_402__flag[0] <= 1'b0;
		ejection_channels_401__flag[0] <= 1'b0;
		ejection_channels_400__flag[0] <= 1'b0;
		ejection_channels_399__flag[0] <= 1'b0;
		ejection_channels_398__flag[0] <= 1'b0;
		ejection_channels_397__flag[0] <= 1'b0;
		ejection_channels_396__flag[0] <= 1'b0;
		ejection_channels_395__flag[0] <= 1'b0;
		ejection_channels_394__flag[0] <= 1'b0;
		ejection_channels_393__flag[0] <= 1'b0;
		ejection_channels_392__flag[0] <= 1'b0;
		ejection_channels_391__flag[0] <= 1'b0;
		ejection_channels_390__flag[0] <= 1'b0;
		ejection_channels_389__flag[0] <= 1'b0;
		ejection_channels_388__flag[0] <= 1'b0;
		ejection_channels_387__flag[0] <= 1'b0;
		ejection_channels_386__flag[0] <= 1'b0;
		ejection_channels_385__flag[0] <= 1'b0;
		ejection_channels_384__flag[0] <= 1'b0;
		ejection_channels_383__flag[0] <= 1'b0;
		ejection_channels_382__flag[0] <= 1'b0;
		ejection_channels_381__flag[0] <= 1'b0;
		ejection_channels_380__flag[0] <= 1'b0;
		ejection_channels_379__flag[0] <= 1'b0;
		ejection_channels_378__flag[0] <= 1'b0;
		ejection_channels_377__flag[0] <= 1'b0;
		ejection_channels_376__flag[0] <= 1'b0;
		ejection_channels_375__flag[0] <= 1'b0;
		ejection_channels_374__flag[0] <= 1'b0;
		ejection_channels_373__flag[0] <= 1'b0;
		ejection_channels_372__flag[0] <= 1'b0;
		ejection_channels_371__flag[0] <= 1'b0;
		ejection_channels_370__flag[0] <= 1'b0;
		ejection_channels_369__flag[0] <= 1'b0;
		ejection_channels_368__flag[0] <= 1'b0;
		ejection_channels_367__flag[0] <= 1'b0;
		ejection_channels_366__flag[0] <= 1'b0;
		ejection_channels_365__flag[0] <= 1'b0;
		ejection_channels_364__flag[0] <= 1'b0;
		ejection_channels_363__flag[0] <= 1'b0;
		ejection_channels_362__flag[0] <= 1'b0;
		ejection_channels_361__flag[0] <= 1'b0;
		ejection_channels_360__flag[0] <= 1'b0;
		ejection_channels_359__flag[0] <= 1'b0;
		ejection_channels_358__flag[0] <= 1'b0;
		ejection_channels_357__flag[0] <= 1'b0;
		ejection_channels_356__flag[0] <= 1'b0;
		ejection_channels_355__flag[0] <= 1'b0;
		ejection_channels_354__flag[0] <= 1'b0;
		ejection_channels_353__flag[0] <= 1'b0;
		ejection_channels_352__flag[0] <= 1'b0;
		ejection_channels_351__flag[0] <= 1'b0;
		ejection_channels_350__flag[0] <= 1'b0;
		ejection_channels_349__flag[0] <= 1'b0;
		ejection_channels_348__flag[0] <= 1'b0;
		ejection_channels_347__flag[0] <= 1'b0;
		ejection_channels_346__flag[0] <= 1'b0;
		ejection_channels_345__flag[0] <= 1'b0;
		ejection_channels_344__flag[0] <= 1'b0;
		ejection_channels_343__flag[0] <= 1'b0;
		ejection_channels_342__flag[0] <= 1'b0;
		ejection_channels_341__flag[0] <= 1'b0;
		ejection_channels_340__flag[0] <= 1'b0;
		ejection_channels_339__flag[0] <= 1'b0;
		ejection_channels_338__flag[0] <= 1'b0;
		ejection_channels_337__flag[0] <= 1'b0;
		ejection_channels_336__flag[0] <= 1'b0;
		ejection_channels_335__flag[0] <= 1'b0;
		ejection_channels_334__flag[0] <= 1'b0;
		ejection_channels_333__flag[0] <= 1'b0;
		ejection_channels_332__flag[0] <= 1'b0;
		ejection_channels_331__flag[0] <= 1'b0;
		ejection_channels_330__flag[0] <= 1'b0;
		ejection_channels_329__flag[0] <= 1'b0;
		ejection_channels_328__flag[0] <= 1'b0;
		ejection_channels_327__flag[0] <= 1'b0;
		ejection_channels_326__flag[0] <= 1'b0;
		ejection_channels_325__flag[0] <= 1'b0;
		ejection_channels_324__flag[0] <= 1'b0;
		ejection_channels_323__flag[0] <= 1'b0;
		ejection_channels_322__flag[0] <= 1'b0;
		ejection_channels_321__flag[0] <= 1'b0;
		ejection_channels_320__flag[0] <= 1'b0;
		ejection_channels_319__flag[0] <= 1'b0;
		ejection_channels_318__flag[0] <= 1'b0;
		ejection_channels_317__flag[0] <= 1'b0;
		ejection_channels_316__flag[0] <= 1'b0;
		ejection_channels_315__flag[0] <= 1'b0;
		ejection_channels_314__flag[0] <= 1'b0;
		ejection_channels_313__flag[0] <= 1'b0;
		ejection_channels_312__flag[0] <= 1'b0;
		ejection_channels_311__flag[0] <= 1'b0;
		ejection_channels_310__flag[0] <= 1'b0;
		ejection_channels_309__flag[0] <= 1'b0;
		ejection_channels_308__flag[0] <= 1'b0;
		ejection_channels_307__flag[0] <= 1'b0;
		ejection_channels_306__flag[0] <= 1'b0;
		ejection_channels_305__flag[0] <= 1'b0;
		ejection_channels_304__flag[0] <= 1'b0;
		ejection_channels_303__flag[0] <= 1'b0;
		ejection_channels_302__flag[0] <= 1'b0;
		ejection_channels_301__flag[0] <= 1'b0;
		ejection_channels_300__flag[0] <= 1'b0;
		ejection_channels_299__flag[0] <= 1'b0;
		ejection_channels_298__flag[0] <= 1'b0;
		ejection_channels_297__flag[0] <= 1'b0;
		ejection_channels_296__flag[0] <= 1'b0;
		ejection_channels_295__flag[0] <= 1'b0;
		ejection_channels_294__flag[0] <= 1'b0;
		ejection_channels_293__flag[0] <= 1'b0;
		ejection_channels_292__flag[0] <= 1'b0;
		ejection_channels_291__flag[0] <= 1'b0;
		ejection_channels_290__flag[0] <= 1'b0;
		ejection_channels_289__flag[0] <= 1'b0;
		ejection_channels_288__flag[0] <= 1'b0;
		ejection_channels_287__flag[0] <= 1'b0;
		ejection_channels_286__flag[0] <= 1'b0;
		ejection_channels_285__flag[0] <= 1'b0;
		ejection_channels_284__flag[0] <= 1'b0;
		ejection_channels_283__flag[0] <= 1'b0;
		ejection_channels_282__flag[0] <= 1'b0;
		ejection_channels_281__flag[0] <= 1'b0;
		ejection_channels_280__flag[0] <= 1'b0;
		ejection_channels_279__flag[0] <= 1'b0;
		ejection_channels_278__flag[0] <= 1'b0;
		ejection_channels_277__flag[0] <= 1'b0;
		ejection_channels_276__flag[0] <= 1'b0;
		ejection_channels_275__flag[0] <= 1'b0;
		ejection_channels_274__flag[0] <= 1'b0;
		ejection_channels_273__flag[0] <= 1'b0;
		ejection_channels_272__flag[0] <= 1'b0;
		ejection_channels_271__flag[0] <= 1'b0;
		ejection_channels_270__flag[0] <= 1'b0;
		ejection_channels_269__flag[0] <= 1'b0;
		ejection_channels_268__flag[0] <= 1'b0;
		ejection_channels_267__flag[0] <= 1'b0;
		ejection_channels_266__flag[0] <= 1'b0;
		ejection_channels_265__flag[0] <= 1'b0;
		ejection_channels_264__flag[0] <= 1'b0;
		ejection_channels_263__flag[0] <= 1'b0;
		ejection_channels_262__flag[0] <= 1'b0;
		ejection_channels_261__flag[0] <= 1'b0;
		ejection_channels_260__flag[0] <= 1'b0;
		ejection_channels_259__flag[0] <= 1'b0;
		ejection_channels_258__flag[0] <= 1'b0;
		ejection_channels_257__flag[0] <= 1'b0;
		ejection_channels_256__flag[0] <= 1'b0;
		ejection_channels_255__flag[0] <= 1'b0;
		ejection_channels_254__flag[0] <= 1'b0;
		ejection_channels_253__flag[0] <= 1'b0;
		ejection_channels_252__flag[0] <= 1'b0;
		ejection_channels_251__flag[0] <= 1'b0;
		ejection_channels_250__flag[0] <= 1'b0;
		ejection_channels_249__flag[0] <= 1'b0;
		ejection_channels_248__flag[0] <= 1'b0;
		ejection_channels_247__flag[0] <= 1'b0;
		ejection_channels_246__flag[0] <= 1'b0;
		ejection_channels_245__flag[0] <= 1'b0;
		ejection_channels_244__flag[0] <= 1'b0;
		ejection_channels_243__flag[0] <= 1'b0;
		ejection_channels_242__flag[0] <= 1'b0;
		ejection_channels_241__flag[0] <= 1'b0;
		ejection_channels_240__flag[0] <= 1'b0;
		ejection_channels_239__flag[0] <= 1'b0;
		ejection_channels_238__flag[0] <= 1'b0;
		ejection_channels_237__flag[0] <= 1'b0;
		ejection_channels_236__flag[0] <= 1'b0;
		ejection_channels_235__flag[0] <= 1'b0;
		ejection_channels_234__flag[0] <= 1'b0;
		ejection_channels_233__flag[0] <= 1'b0;
		ejection_channels_232__flag[0] <= 1'b0;
		ejection_channels_231__flag[0] <= 1'b0;
		ejection_channels_230__flag[0] <= 1'b0;
		ejection_channels_229__flag[0] <= 1'b0;
		ejection_channels_228__flag[0] <= 1'b0;
		ejection_channels_227__flag[0] <= 1'b0;
		ejection_channels_226__flag[0] <= 1'b0;
		ejection_channels_225__flag[0] <= 1'b0;
		ejection_channels_224__flag[0] <= 1'b0;
		ejection_channels_223__flag[0] <= 1'b0;
		ejection_channels_222__flag[0] <= 1'b0;
		ejection_channels_221__flag[0] <= 1'b0;
		ejection_channels_220__flag[0] <= 1'b0;
		ejection_channels_219__flag[0] <= 1'b0;
		ejection_channels_218__flag[0] <= 1'b0;
		ejection_channels_217__flag[0] <= 1'b0;
		ejection_channels_216__flag[0] <= 1'b0;
		ejection_channels_215__flag[0] <= 1'b0;
		ejection_channels_214__flag[0] <= 1'b0;
		ejection_channels_213__flag[0] <= 1'b0;
		ejection_channels_212__flag[0] <= 1'b0;
		ejection_channels_211__flag[0] <= 1'b0;
		ejection_channels_210__flag[0] <= 1'b0;
		ejection_channels_209__flag[0] <= 1'b0;
		ejection_channels_208__flag[0] <= 1'b0;
		ejection_channels_207__flag[0] <= 1'b0;
		ejection_channels_206__flag[0] <= 1'b0;
		ejection_channels_205__flag[0] <= 1'b0;
		ejection_channels_204__flag[0] <= 1'b0;
		ejection_channels_203__flag[0] <= 1'b0;
		ejection_channels_202__flag[0] <= 1'b0;
		ejection_channels_201__flag[0] <= 1'b0;
		ejection_channels_200__flag[0] <= 1'b0;
		ejection_channels_199__flag[0] <= 1'b0;
		ejection_channels_198__flag[0] <= 1'b0;
		ejection_channels_197__flag[0] <= 1'b0;
		ejection_channels_196__flag[0] <= 1'b0;
		ejection_channels_195__flag[0] <= 1'b0;
		ejection_channels_194__flag[0] <= 1'b0;
		ejection_channels_193__flag[0] <= 1'b0;
		ejection_channels_192__flag[0] <= 1'b0;
		ejection_channels_191__flag[0] <= 1'b0;
		ejection_channels_190__flag[0] <= 1'b0;
		ejection_channels_189__flag[0] <= 1'b0;
		ejection_channels_188__flag[0] <= 1'b0;
		ejection_channels_187__flag[0] <= 1'b0;
		ejection_channels_186__flag[0] <= 1'b0;
		ejection_channels_185__flag[0] <= 1'b0;
		ejection_channels_184__flag[0] <= 1'b0;
		ejection_channels_183__flag[0] <= 1'b0;
		ejection_channels_182__flag[0] <= 1'b0;
		ejection_channels_181__flag[0] <= 1'b0;
		ejection_channels_180__flag[0] <= 1'b0;
		ejection_channels_179__flag[0] <= 1'b0;
		ejection_channels_178__flag[0] <= 1'b0;
		ejection_channels_177__flag[0] <= 1'b0;
		ejection_channels_176__flag[0] <= 1'b0;
		ejection_channels_175__flag[0] <= 1'b0;
		ejection_channels_174__flag[0] <= 1'b0;
		ejection_channels_173__flag[0] <= 1'b0;
		ejection_channels_172__flag[0] <= 1'b0;
		ejection_channels_171__flag[0] <= 1'b0;
		ejection_channels_170__flag[0] <= 1'b0;
		ejection_channels_169__flag[0] <= 1'b0;
		ejection_channels_168__flag[0] <= 1'b0;
		ejection_channels_167__flag[0] <= 1'b0;
		ejection_channels_166__flag[0] <= 1'b0;
		ejection_channels_165__flag[0] <= 1'b0;
		ejection_channels_164__flag[0] <= 1'b0;
		ejection_channels_163__flag[0] <= 1'b0;
		ejection_channels_162__flag[0] <= 1'b0;
		ejection_channels_161__flag[0] <= 1'b0;
		ejection_channels_160__flag[0] <= 1'b0;
		ejection_channels_159__flag[0] <= 1'b0;
		ejection_channels_158__flag[0] <= 1'b0;
		ejection_channels_157__flag[0] <= 1'b0;
		ejection_channels_156__flag[0] <= 1'b0;
		ejection_channels_155__flag[0] <= 1'b0;
		ejection_channels_154__flag[0] <= 1'b0;
		ejection_channels_153__flag[0] <= 1'b0;
		ejection_channels_152__flag[0] <= 1'b0;
		ejection_channels_151__flag[0] <= 1'b0;
		ejection_channels_150__flag[0] <= 1'b0;
		ejection_channels_149__flag[0] <= 1'b0;
		ejection_channels_148__flag[0] <= 1'b0;
		ejection_channels_147__flag[0] <= 1'b0;
		ejection_channels_146__flag[0] <= 1'b0;
		ejection_channels_145__flag[0] <= 1'b0;
		ejection_channels_144__flag[0] <= 1'b0;
		ejection_channels_143__flag[0] <= 1'b0;
		ejection_channels_142__flag[0] <= 1'b0;
		ejection_channels_141__flag[0] <= 1'b0;
		ejection_channels_140__flag[0] <= 1'b0;
		ejection_channels_139__flag[0] <= 1'b0;
		ejection_channels_138__flag[0] <= 1'b0;
		ejection_channels_137__flag[0] <= 1'b0;
		ejection_channels_136__flag[0] <= 1'b0;
		ejection_channels_135__flag[0] <= 1'b0;
		ejection_channels_134__flag[0] <= 1'b0;
		ejection_channels_133__flag[0] <= 1'b0;
		ejection_channels_132__flag[0] <= 1'b0;
		ejection_channels_131__flag[0] <= 1'b0;
		ejection_channels_130__flag[0] <= 1'b0;
		ejection_channels_129__flag[0] <= 1'b0;
		ejection_channels_128__flag[0] <= 1'b0;
		ejection_channels_127__flag[0] <= 1'b0;
		ejection_channels_126__flag[0] <= 1'b0;
		ejection_channels_125__flag[0] <= 1'b0;
		ejection_channels_124__flag[0] <= 1'b0;
		ejection_channels_123__flag[0] <= 1'b0;
		ejection_channels_122__flag[0] <= 1'b0;
		ejection_channels_121__flag[0] <= 1'b0;
		ejection_channels_120__flag[0] <= 1'b0;
		ejection_channels_119__flag[0] <= 1'b0;
		ejection_channels_118__flag[0] <= 1'b0;
		ejection_channels_117__flag[0] <= 1'b0;
		ejection_channels_116__flag[0] <= 1'b0;
		ejection_channels_115__flag[0] <= 1'b0;
		ejection_channels_114__flag[0] <= 1'b0;
		ejection_channels_113__flag[0] <= 1'b0;
		ejection_channels_112__flag[0] <= 1'b0;
		ejection_channels_111__flag[0] <= 1'b0;
		ejection_channels_110__flag[0] <= 1'b0;
		ejection_channels_109__flag[0] <= 1'b0;
		ejection_channels_108__flag[0] <= 1'b0;
		ejection_channels_107__flag[0] <= 1'b0;
		ejection_channels_106__flag[0] <= 1'b0;
		ejection_channels_105__flag[0] <= 1'b0;
		ejection_channels_104__flag[0] <= 1'b0;
		ejection_channels_103__flag[0] <= 1'b0;
		ejection_channels_102__flag[0] <= 1'b0;
		ejection_channels_101__flag[0] <= 1'b0;
		ejection_channels_100__flag[0] <= 1'b0;
		ejection_channels_99__flag[0] <= 1'b0;
		ejection_channels_98__flag[0] <= 1'b0;
		ejection_channels_97__flag[0] <= 1'b0;
		ejection_channels_96__flag[0] <= 1'b0;
		ejection_channels_95__flag[0] <= 1'b0;
		ejection_channels_94__flag[0] <= 1'b0;
		ejection_channels_93__flag[0] <= 1'b0;
		ejection_channels_92__flag[0] <= 1'b0;
		ejection_channels_91__flag[0] <= 1'b0;
		ejection_channels_90__flag[0] <= 1'b0;
		ejection_channels_89__flag[0] <= 1'b0;
		ejection_channels_88__flag[0] <= 1'b0;
		ejection_channels_87__flag[0] <= 1'b0;
		ejection_channels_86__flag[0] <= 1'b0;
		ejection_channels_85__flag[0] <= 1'b0;
		ejection_channels_84__flag[0] <= 1'b0;
		ejection_channels_83__flag[0] <= 1'b0;
		ejection_channels_82__flag[0] <= 1'b0;
		ejection_channels_81__flag[0] <= 1'b0;
		ejection_channels_80__flag[0] <= 1'b0;
		ejection_channels_79__flag[0] <= 1'b0;
		ejection_channels_78__flag[0] <= 1'b0;
		ejection_channels_77__flag[0] <= 1'b0;
		ejection_channels_76__flag[0] <= 1'b0;
		ejection_channels_75__flag[0] <= 1'b0;
		ejection_channels_74__flag[0] <= 1'b0;
		ejection_channels_73__flag[0] <= 1'b0;
		ejection_channels_72__flag[0] <= 1'b0;
		ejection_channels_71__flag[0] <= 1'b0;
		ejection_channels_70__flag[0] <= 1'b0;
		ejection_channels_69__flag[0] <= 1'b0;
		ejection_channels_68__flag[0] <= 1'b0;
		ejection_channels_67__flag[0] <= 1'b0;
		ejection_channels_66__flag[0] <= 1'b0;
		ejection_channels_65__flag[0] <= 1'b0;
		ejection_channels_64__flag[0] <= 1'b0;
		ejection_channels_63__flag[0] <= 1'b0;
		ejection_channels_62__flag[0] <= 1'b0;
		ejection_channels_61__flag[0] <= 1'b0;
		ejection_channels_60__flag[0] <= 1'b0;
		ejection_channels_59__flag[0] <= 1'b0;
		ejection_channels_58__flag[0] <= 1'b0;
		ejection_channels_57__flag[0] <= 1'b0;
		ejection_channels_56__flag[0] <= 1'b0;
		ejection_channels_55__flag[0] <= 1'b0;
		ejection_channels_54__flag[0] <= 1'b0;
		ejection_channels_53__flag[0] <= 1'b0;
		ejection_channels_52__flag[0] <= 1'b0;
		ejection_channels_51__flag[0] <= 1'b0;
		ejection_channels_50__flag[0] <= 1'b0;
		ejection_channels_49__flag[0] <= 1'b0;
		ejection_channels_48__flag[0] <= 1'b0;
		ejection_channels_47__flag[0] <= 1'b0;
		ejection_channels_46__flag[0] <= 1'b0;
		ejection_channels_45__flag[0] <= 1'b0;
		ejection_channels_44__flag[0] <= 1'b0;
		ejection_channels_43__flag[0] <= 1'b0;
		ejection_channels_42__flag[0] <= 1'b0;
		ejection_channels_41__flag[0] <= 1'b0;
		ejection_channels_40__flag[0] <= 1'b0;
		ejection_channels_39__flag[0] <= 1'b0;
		ejection_channels_38__flag[0] <= 1'b0;
		ejection_channels_37__flag[0] <= 1'b0;
		ejection_channels_36__flag[0] <= 1'b0;
		ejection_channels_35__flag[0] <= 1'b0;
		ejection_channels_34__flag[0] <= 1'b0;
		ejection_channels_33__flag[0] <= 1'b0;
		ejection_channels_32__flag[0] <= 1'b0;
		ejection_channels_31__flag[0] <= 1'b0;
		ejection_channels_30__flag[0] <= 1'b0;
		ejection_channels_29__flag[0] <= 1'b0;
		ejection_channels_28__flag[0] <= 1'b0;
		ejection_channels_27__flag[0] <= 1'b0;
		ejection_channels_26__flag[0] <= 1'b0;
		ejection_channels_25__flag[0] <= 1'b0;
		ejection_channels_24__flag[0] <= 1'b0;
		ejection_channels_23__flag[0] <= 1'b0;
		ejection_channels_22__flag[0] <= 1'b0;
		ejection_channels_21__flag[0] <= 1'b0;
		ejection_channels_20__flag[0] <= 1'b0;
		ejection_channels_19__flag[0] <= 1'b0;
		ejection_channels_18__flag[0] <= 1'b0;
		ejection_channels_17__flag[0] <= 1'b0;
		ejection_channels_16__flag[0] <= 1'b0;
		ejection_channels_15__flag[0] <= 1'b0;
		ejection_channels_14__flag[0] <= 1'b0;
		ejection_channels_13__flag[0] <= 1'b0;
		ejection_channels_12__flag[0] <= 1'b0;
		ejection_channels_11__flag[0] <= 1'b0;
		ejection_channels_10__flag[0] <= 1'b0;
		ejection_channels_9__flag[0] <= 1'b0;
		ejection_channels_8__flag[0] <= 1'b0;
		ejection_channels_7__flag[0] <= 1'b0;
		ejection_channels_6__flag[0] <= 1'b0;
		ejection_channels_5__flag[0] <= 1'b0;
		ejection_channels_4__flag[0] <= 1'b0;
		ejection_channels_3__flag[0] <= 1'b0;
		ejection_channels_2__flag[0] <= 1'b0;
		ejection_channels_1__flag[0] <= 1'b0;
		ejection_channels_0__flag[0] <= 1'b0;
		rtr_error_8__flag[0] <= 1'b0;
		rtr_error_7__flag[0] <= 1'b0;
		rtr_error_6__flag[0] <= 1'b0;
		rtr_error_5__flag[0] <= 1'b0;
		rtr_error_4__flag[0] <= 1'b0;
		rtr_error_3__flag[0] <= 1'b0;
		rtr_error_2__flag[0] <= 1'b0;
		rtr_error_1__flag[0] <= 1'b0;
		rtr_error_0__flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge clk[0]) begin
		reset <= $random;
		injection_channels_629_ <= $random;
		injection_channels_628_ <= $random;
		injection_channels_627_ <= $random;
		injection_channels_626_ <= $random;
		injection_channels_625_ <= $random;
		injection_channels_624_ <= $random;
		injection_channels_623_ <= $random;
		injection_channels_622_ <= $random;
		injection_channels_621_ <= $random;
		injection_channels_620_ <= $random;
		injection_channels_619_ <= $random;
		injection_channels_618_ <= $random;
		injection_channels_617_ <= $random;
		injection_channels_616_ <= $random;
		injection_channels_615_ <= $random;
		injection_channels_614_ <= $random;
		injection_channels_613_ <= $random;
		injection_channels_612_ <= $random;
		injection_channels_611_ <= $random;
		injection_channels_610_ <= $random;
		injection_channels_609_ <= $random;
		injection_channels_608_ <= $random;
		injection_channels_607_ <= $random;
		injection_channels_606_ <= $random;
		injection_channels_605_ <= $random;
		injection_channels_604_ <= $random;
		injection_channels_603_ <= $random;
		injection_channels_602_ <= $random;
		injection_channels_601_ <= $random;
		injection_channels_600_ <= $random;
		injection_channels_599_ <= $random;
		injection_channels_598_ <= $random;
		injection_channels_597_ <= $random;
		injection_channels_596_ <= $random;
		injection_channels_595_ <= $random;
		injection_channels_594_ <= $random;
		injection_channels_593_ <= $random;
		injection_channels_592_ <= $random;
		injection_channels_591_ <= $random;
		injection_channels_590_ <= $random;
		injection_channels_589_ <= $random;
		injection_channels_588_ <= $random;
		injection_channels_587_ <= $random;
		injection_channels_586_ <= $random;
		injection_channels_585_ <= $random;
		injection_channels_584_ <= $random;
		injection_channels_583_ <= $random;
		injection_channels_582_ <= $random;
		injection_channels_581_ <= $random;
		injection_channels_580_ <= $random;
		injection_channels_579_ <= $random;
		injection_channels_578_ <= $random;
		injection_channels_577_ <= $random;
		injection_channels_576_ <= $random;
		injection_channels_575_ <= $random;
		injection_channels_574_ <= $random;
		injection_channels_573_ <= $random;
		injection_channels_572_ <= $random;
		injection_channels_571_ <= $random;
		injection_channels_570_ <= $random;
		injection_channels_569_ <= $random;
		injection_channels_568_ <= $random;
		injection_channels_567_ <= $random;
		injection_channels_566_ <= $random;
		injection_channels_565_ <= $random;
		injection_channels_564_ <= $random;
		injection_channels_563_ <= $random;
		injection_channels_562_ <= $random;
		injection_channels_561_ <= $random;
		injection_channels_560_ <= $random;
		injection_channels_559_ <= $random;
		injection_channels_558_ <= $random;
		injection_channels_557_ <= $random;
		injection_channels_556_ <= $random;
		injection_channels_555_ <= $random;
		injection_channels_554_ <= $random;
		injection_channels_553_ <= $random;
		injection_channels_552_ <= $random;
		injection_channels_551_ <= $random;
		injection_channels_550_ <= $random;
		injection_channels_549_ <= $random;
		injection_channels_548_ <= $random;
		injection_channels_547_ <= $random;
		injection_channels_546_ <= $random;
		injection_channels_545_ <= $random;
		injection_channels_544_ <= $random;
		injection_channels_543_ <= $random;
		injection_channels_542_ <= $random;
		injection_channels_541_ <= $random;
		injection_channels_540_ <= $random;
		injection_channels_539_ <= $random;
		injection_channels_538_ <= $random;
		injection_channels_537_ <= $random;
		injection_channels_536_ <= $random;
		injection_channels_535_ <= $random;
		injection_channels_534_ <= $random;
		injection_channels_533_ <= $random;
		injection_channels_532_ <= $random;
		injection_channels_531_ <= $random;
		injection_channels_530_ <= $random;
		injection_channels_529_ <= $random;
		injection_channels_528_ <= $random;
		injection_channels_527_ <= $random;
		injection_channels_526_ <= $random;
		injection_channels_525_ <= $random;
		injection_channels_524_ <= $random;
		injection_channels_523_ <= $random;
		injection_channels_522_ <= $random;
		injection_channels_521_ <= $random;
		injection_channels_520_ <= $random;
		injection_channels_519_ <= $random;
		injection_channels_518_ <= $random;
		injection_channels_517_ <= $random;
		injection_channels_516_ <= $random;
		injection_channels_515_ <= $random;
		injection_channels_514_ <= $random;
		injection_channels_513_ <= $random;
		injection_channels_512_ <= $random;
		injection_channels_511_ <= $random;
		injection_channels_510_ <= $random;
		injection_channels_509_ <= $random;
		injection_channels_508_ <= $random;
		injection_channels_507_ <= $random;
		injection_channels_506_ <= $random;
		injection_channels_505_ <= $random;
		injection_channels_504_ <= $random;
		injection_channels_503_ <= $random;
		injection_channels_502_ <= $random;
		injection_channels_501_ <= $random;
		injection_channels_500_ <= $random;
		injection_channels_499_ <= $random;
		injection_channels_498_ <= $random;
		injection_channels_497_ <= $random;
		injection_channels_496_ <= $random;
		injection_channels_495_ <= $random;
		injection_channels_494_ <= $random;
		injection_channels_493_ <= $random;
		injection_channels_492_ <= $random;
		injection_channels_491_ <= $random;
		injection_channels_490_ <= $random;
		injection_channels_489_ <= $random;
		injection_channels_488_ <= $random;
		injection_channels_487_ <= $random;
		injection_channels_486_ <= $random;
		injection_channels_485_ <= $random;
		injection_channels_484_ <= $random;
		injection_channels_483_ <= $random;
		injection_channels_482_ <= $random;
		injection_channels_481_ <= $random;
		injection_channels_480_ <= $random;
		injection_channels_479_ <= $random;
		injection_channels_478_ <= $random;
		injection_channels_477_ <= $random;
		injection_channels_476_ <= $random;
		injection_channels_475_ <= $random;
		injection_channels_474_ <= $random;
		injection_channels_473_ <= $random;
		injection_channels_472_ <= $random;
		injection_channels_471_ <= $random;
		injection_channels_470_ <= $random;
		injection_channels_469_ <= $random;
		injection_channels_468_ <= $random;
		injection_channels_467_ <= $random;
		injection_channels_466_ <= $random;
		injection_channels_465_ <= $random;
		injection_channels_464_ <= $random;
		injection_channels_463_ <= $random;
		injection_channels_462_ <= $random;
		injection_channels_461_ <= $random;
		injection_channels_460_ <= $random;
		injection_channels_459_ <= $random;
		injection_channels_458_ <= $random;
		injection_channels_457_ <= $random;
		injection_channels_456_ <= $random;
		injection_channels_455_ <= $random;
		injection_channels_454_ <= $random;
		injection_channels_453_ <= $random;
		injection_channels_452_ <= $random;
		injection_channels_451_ <= $random;
		injection_channels_450_ <= $random;
		injection_channels_449_ <= $random;
		injection_channels_448_ <= $random;
		injection_channels_447_ <= $random;
		injection_channels_446_ <= $random;
		injection_channels_445_ <= $random;
		injection_channels_444_ <= $random;
		injection_channels_443_ <= $random;
		injection_channels_442_ <= $random;
		injection_channels_441_ <= $random;
		injection_channels_440_ <= $random;
		injection_channels_439_ <= $random;
		injection_channels_438_ <= $random;
		injection_channels_437_ <= $random;
		injection_channels_436_ <= $random;
		injection_channels_435_ <= $random;
		injection_channels_434_ <= $random;
		injection_channels_433_ <= $random;
		injection_channels_432_ <= $random;
		injection_channels_431_ <= $random;
		injection_channels_430_ <= $random;
		injection_channels_429_ <= $random;
		injection_channels_428_ <= $random;
		injection_channels_427_ <= $random;
		injection_channels_426_ <= $random;
		injection_channels_425_ <= $random;
		injection_channels_424_ <= $random;
		injection_channels_423_ <= $random;
		injection_channels_422_ <= $random;
		injection_channels_421_ <= $random;
		injection_channels_420_ <= $random;
		injection_channels_419_ <= $random;
		injection_channels_418_ <= $random;
		injection_channels_417_ <= $random;
		injection_channels_416_ <= $random;
		injection_channels_415_ <= $random;
		injection_channels_414_ <= $random;
		injection_channels_413_ <= $random;
		injection_channels_412_ <= $random;
		injection_channels_411_ <= $random;
		injection_channels_410_ <= $random;
		injection_channels_409_ <= $random;
		injection_channels_408_ <= $random;
		injection_channels_407_ <= $random;
		injection_channels_406_ <= $random;
		injection_channels_405_ <= $random;
		injection_channels_404_ <= $random;
		injection_channels_403_ <= $random;
		injection_channels_402_ <= $random;
		injection_channels_401_ <= $random;
		injection_channels_400_ <= $random;
		injection_channels_399_ <= $random;
		injection_channels_398_ <= $random;
		injection_channels_397_ <= $random;
		injection_channels_396_ <= $random;
		injection_channels_395_ <= $random;
		injection_channels_394_ <= $random;
		injection_channels_393_ <= $random;
		injection_channels_392_ <= $random;
		injection_channels_391_ <= $random;
		injection_channels_390_ <= $random;
		injection_channels_389_ <= $random;
		injection_channels_388_ <= $random;
		injection_channels_387_ <= $random;
		injection_channels_386_ <= $random;
		injection_channels_385_ <= $random;
		injection_channels_384_ <= $random;
		injection_channels_383_ <= $random;
		injection_channels_382_ <= $random;
		injection_channels_381_ <= $random;
		injection_channels_380_ <= $random;
		injection_channels_379_ <= $random;
		injection_channels_378_ <= $random;
		injection_channels_377_ <= $random;
		injection_channels_376_ <= $random;
		injection_channels_375_ <= $random;
		injection_channels_374_ <= $random;
		injection_channels_373_ <= $random;
		injection_channels_372_ <= $random;
		injection_channels_371_ <= $random;
		injection_channels_370_ <= $random;
		injection_channels_369_ <= $random;
		injection_channels_368_ <= $random;
		injection_channels_367_ <= $random;
		injection_channels_366_ <= $random;
		injection_channels_365_ <= $random;
		injection_channels_364_ <= $random;
		injection_channels_363_ <= $random;
		injection_channels_362_ <= $random;
		injection_channels_361_ <= $random;
		injection_channels_360_ <= $random;
		injection_channels_359_ <= $random;
		injection_channels_358_ <= $random;
		injection_channels_357_ <= $random;
		injection_channels_356_ <= $random;
		injection_channels_355_ <= $random;
		injection_channels_354_ <= $random;
		injection_channels_353_ <= $random;
		injection_channels_352_ <= $random;
		injection_channels_351_ <= $random;
		injection_channels_350_ <= $random;
		injection_channels_349_ <= $random;
		injection_channels_348_ <= $random;
		injection_channels_347_ <= $random;
		injection_channels_346_ <= $random;
		injection_channels_345_ <= $random;
		injection_channels_344_ <= $random;
		injection_channels_343_ <= $random;
		injection_channels_342_ <= $random;
		injection_channels_341_ <= $random;
		injection_channels_340_ <= $random;
		injection_channels_339_ <= $random;
		injection_channels_338_ <= $random;
		injection_channels_337_ <= $random;
		injection_channels_336_ <= $random;
		injection_channels_335_ <= $random;
		injection_channels_334_ <= $random;
		injection_channels_333_ <= $random;
		injection_channels_332_ <= $random;
		injection_channels_331_ <= $random;
		injection_channels_330_ <= $random;
		injection_channels_329_ <= $random;
		injection_channels_328_ <= $random;
		injection_channels_327_ <= $random;
		injection_channels_326_ <= $random;
		injection_channels_325_ <= $random;
		injection_channels_324_ <= $random;
		injection_channels_323_ <= $random;
		injection_channels_322_ <= $random;
		injection_channels_321_ <= $random;
		injection_channels_320_ <= $random;
		injection_channels_319_ <= $random;
		injection_channels_318_ <= $random;
		injection_channels_317_ <= $random;
		injection_channels_316_ <= $random;
		injection_channels_315_ <= $random;
		injection_channels_314_ <= $random;
		injection_channels_313_ <= $random;
		injection_channels_312_ <= $random;
		injection_channels_311_ <= $random;
		injection_channels_310_ <= $random;
		injection_channels_309_ <= $random;
		injection_channels_308_ <= $random;
		injection_channels_307_ <= $random;
		injection_channels_306_ <= $random;
		injection_channels_305_ <= $random;
		injection_channels_304_ <= $random;
		injection_channels_303_ <= $random;
		injection_channels_302_ <= $random;
		injection_channels_301_ <= $random;
		injection_channels_300_ <= $random;
		injection_channels_299_ <= $random;
		injection_channels_298_ <= $random;
		injection_channels_297_ <= $random;
		injection_channels_296_ <= $random;
		injection_channels_295_ <= $random;
		injection_channels_294_ <= $random;
		injection_channels_293_ <= $random;
		injection_channels_292_ <= $random;
		injection_channels_291_ <= $random;
		injection_channels_290_ <= $random;
		injection_channels_289_ <= $random;
		injection_channels_288_ <= $random;
		injection_channels_287_ <= $random;
		injection_channels_286_ <= $random;
		injection_channels_285_ <= $random;
		injection_channels_284_ <= $random;
		injection_channels_283_ <= $random;
		injection_channels_282_ <= $random;
		injection_channels_281_ <= $random;
		injection_channels_280_ <= $random;
		injection_channels_279_ <= $random;
		injection_channels_278_ <= $random;
		injection_channels_277_ <= $random;
		injection_channels_276_ <= $random;
		injection_channels_275_ <= $random;
		injection_channels_274_ <= $random;
		injection_channels_273_ <= $random;
		injection_channels_272_ <= $random;
		injection_channels_271_ <= $random;
		injection_channels_270_ <= $random;
		injection_channels_269_ <= $random;
		injection_channels_268_ <= $random;
		injection_channels_267_ <= $random;
		injection_channels_266_ <= $random;
		injection_channels_265_ <= $random;
		injection_channels_264_ <= $random;
		injection_channels_263_ <= $random;
		injection_channels_262_ <= $random;
		injection_channels_261_ <= $random;
		injection_channels_260_ <= $random;
		injection_channels_259_ <= $random;
		injection_channels_258_ <= $random;
		injection_channels_257_ <= $random;
		injection_channels_256_ <= $random;
		injection_channels_255_ <= $random;
		injection_channels_254_ <= $random;
		injection_channels_253_ <= $random;
		injection_channels_252_ <= $random;
		injection_channels_251_ <= $random;
		injection_channels_250_ <= $random;
		injection_channels_249_ <= $random;
		injection_channels_248_ <= $random;
		injection_channels_247_ <= $random;
		injection_channels_246_ <= $random;
		injection_channels_245_ <= $random;
		injection_channels_244_ <= $random;
		injection_channels_243_ <= $random;
		injection_channels_242_ <= $random;
		injection_channels_241_ <= $random;
		injection_channels_240_ <= $random;
		injection_channels_239_ <= $random;
		injection_channels_238_ <= $random;
		injection_channels_237_ <= $random;
		injection_channels_236_ <= $random;
		injection_channels_235_ <= $random;
		injection_channels_234_ <= $random;
		injection_channels_233_ <= $random;
		injection_channels_232_ <= $random;
		injection_channels_231_ <= $random;
		injection_channels_230_ <= $random;
		injection_channels_229_ <= $random;
		injection_channels_228_ <= $random;
		injection_channels_227_ <= $random;
		injection_channels_226_ <= $random;
		injection_channels_225_ <= $random;
		injection_channels_224_ <= $random;
		injection_channels_223_ <= $random;
		injection_channels_222_ <= $random;
		injection_channels_221_ <= $random;
		injection_channels_220_ <= $random;
		injection_channels_219_ <= $random;
		injection_channels_218_ <= $random;
		injection_channels_217_ <= $random;
		injection_channels_216_ <= $random;
		injection_channels_215_ <= $random;
		injection_channels_214_ <= $random;
		injection_channels_213_ <= $random;
		injection_channels_212_ <= $random;
		injection_channels_211_ <= $random;
		injection_channels_210_ <= $random;
		injection_channels_209_ <= $random;
		injection_channels_208_ <= $random;
		injection_channels_207_ <= $random;
		injection_channels_206_ <= $random;
		injection_channels_205_ <= $random;
		injection_channels_204_ <= $random;
		injection_channels_203_ <= $random;
		injection_channels_202_ <= $random;
		injection_channels_201_ <= $random;
		injection_channels_200_ <= $random;
		injection_channels_199_ <= $random;
		injection_channels_198_ <= $random;
		injection_channels_197_ <= $random;
		injection_channels_196_ <= $random;
		injection_channels_195_ <= $random;
		injection_channels_194_ <= $random;
		injection_channels_193_ <= $random;
		injection_channels_192_ <= $random;
		injection_channels_191_ <= $random;
		injection_channels_190_ <= $random;
		injection_channels_189_ <= $random;
		injection_channels_188_ <= $random;
		injection_channels_187_ <= $random;
		injection_channels_186_ <= $random;
		injection_channels_185_ <= $random;
		injection_channels_184_ <= $random;
		injection_channels_183_ <= $random;
		injection_channels_182_ <= $random;
		injection_channels_181_ <= $random;
		injection_channels_180_ <= $random;
		injection_channels_179_ <= $random;
		injection_channels_178_ <= $random;
		injection_channels_177_ <= $random;
		injection_channels_176_ <= $random;
		injection_channels_175_ <= $random;
		injection_channels_174_ <= $random;
		injection_channels_173_ <= $random;
		injection_channels_172_ <= $random;
		injection_channels_171_ <= $random;
		injection_channels_170_ <= $random;
		injection_channels_169_ <= $random;
		injection_channels_168_ <= $random;
		injection_channels_167_ <= $random;
		injection_channels_166_ <= $random;
		injection_channels_165_ <= $random;
		injection_channels_164_ <= $random;
		injection_channels_163_ <= $random;
		injection_channels_162_ <= $random;
		injection_channels_161_ <= $random;
		injection_channels_160_ <= $random;
		injection_channels_159_ <= $random;
		injection_channels_158_ <= $random;
		injection_channels_157_ <= $random;
		injection_channels_156_ <= $random;
		injection_channels_155_ <= $random;
		injection_channels_154_ <= $random;
		injection_channels_153_ <= $random;
		injection_channels_152_ <= $random;
		injection_channels_151_ <= $random;
		injection_channels_150_ <= $random;
		injection_channels_149_ <= $random;
		injection_channels_148_ <= $random;
		injection_channels_147_ <= $random;
		injection_channels_146_ <= $random;
		injection_channels_145_ <= $random;
		injection_channels_144_ <= $random;
		injection_channels_143_ <= $random;
		injection_channels_142_ <= $random;
		injection_channels_141_ <= $random;
		injection_channels_140_ <= $random;
		injection_channels_139_ <= $random;
		injection_channels_138_ <= $random;
		injection_channels_137_ <= $random;
		injection_channels_136_ <= $random;
		injection_channels_135_ <= $random;
		injection_channels_134_ <= $random;
		injection_channels_133_ <= $random;
		injection_channels_132_ <= $random;
		injection_channels_131_ <= $random;
		injection_channels_130_ <= $random;
		injection_channels_129_ <= $random;
		injection_channels_128_ <= $random;
		injection_channels_127_ <= $random;
		injection_channels_126_ <= $random;
		injection_channels_125_ <= $random;
		injection_channels_124_ <= $random;
		injection_channels_123_ <= $random;
		injection_channels_122_ <= $random;
		injection_channels_121_ <= $random;
		injection_channels_120_ <= $random;
		injection_channels_119_ <= $random;
		injection_channels_118_ <= $random;
		injection_channels_117_ <= $random;
		injection_channels_116_ <= $random;
		injection_channels_115_ <= $random;
		injection_channels_114_ <= $random;
		injection_channels_113_ <= $random;
		injection_channels_112_ <= $random;
		injection_channels_111_ <= $random;
		injection_channels_110_ <= $random;
		injection_channels_109_ <= $random;
		injection_channels_108_ <= $random;
		injection_channels_107_ <= $random;
		injection_channels_106_ <= $random;
		injection_channels_105_ <= $random;
		injection_channels_104_ <= $random;
		injection_channels_103_ <= $random;
		injection_channels_102_ <= $random;
		injection_channels_101_ <= $random;
		injection_channels_100_ <= $random;
		injection_channels_99_ <= $random;
		injection_channels_98_ <= $random;
		injection_channels_97_ <= $random;
		injection_channels_96_ <= $random;
		injection_channels_95_ <= $random;
		injection_channels_94_ <= $random;
		injection_channels_93_ <= $random;
		injection_channels_92_ <= $random;
		injection_channels_91_ <= $random;
		injection_channels_90_ <= $random;
		injection_channels_89_ <= $random;
		injection_channels_88_ <= $random;
		injection_channels_87_ <= $random;
		injection_channels_86_ <= $random;
		injection_channels_85_ <= $random;
		injection_channels_84_ <= $random;
		injection_channels_83_ <= $random;
		injection_channels_82_ <= $random;
		injection_channels_81_ <= $random;
		injection_channels_80_ <= $random;
		injection_channels_79_ <= $random;
		injection_channels_78_ <= $random;
		injection_channels_77_ <= $random;
		injection_channels_76_ <= $random;
		injection_channels_75_ <= $random;
		injection_channels_74_ <= $random;
		injection_channels_73_ <= $random;
		injection_channels_72_ <= $random;
		injection_channels_71_ <= $random;
		injection_channels_70_ <= $random;
		injection_channels_69_ <= $random;
		injection_channels_68_ <= $random;
		injection_channels_67_ <= $random;
		injection_channels_66_ <= $random;
		injection_channels_65_ <= $random;
		injection_channels_64_ <= $random;
		injection_channels_63_ <= $random;
		injection_channels_62_ <= $random;
		injection_channels_61_ <= $random;
		injection_channels_60_ <= $random;
		injection_channels_59_ <= $random;
		injection_channels_58_ <= $random;
		injection_channels_57_ <= $random;
		injection_channels_56_ <= $random;
		injection_channels_55_ <= $random;
		injection_channels_54_ <= $random;
		injection_channels_53_ <= $random;
		injection_channels_52_ <= $random;
		injection_channels_51_ <= $random;
		injection_channels_50_ <= $random;
		injection_channels_49_ <= $random;
		injection_channels_48_ <= $random;
		injection_channels_47_ <= $random;
		injection_channels_46_ <= $random;
		injection_channels_45_ <= $random;
		injection_channels_44_ <= $random;
		injection_channels_43_ <= $random;
		injection_channels_42_ <= $random;
		injection_channels_41_ <= $random;
		injection_channels_40_ <= $random;
		injection_channels_39_ <= $random;
		injection_channels_38_ <= $random;
		injection_channels_37_ <= $random;
		injection_channels_36_ <= $random;
		injection_channels_35_ <= $random;
		injection_channels_34_ <= $random;
		injection_channels_33_ <= $random;
		injection_channels_32_ <= $random;
		injection_channels_31_ <= $random;
		injection_channels_30_ <= $random;
		injection_channels_29_ <= $random;
		injection_channels_28_ <= $random;
		injection_channels_27_ <= $random;
		injection_channels_26_ <= $random;
		injection_channels_25_ <= $random;
		injection_channels_24_ <= $random;
		injection_channels_23_ <= $random;
		injection_channels_22_ <= $random;
		injection_channels_21_ <= $random;
		injection_channels_20_ <= $random;
		injection_channels_19_ <= $random;
		injection_channels_18_ <= $random;
		injection_channels_17_ <= $random;
		injection_channels_16_ <= $random;
		injection_channels_15_ <= $random;
		injection_channels_14_ <= $random;
		injection_channels_13_ <= $random;
		injection_channels_12_ <= $random;
		injection_channels_11_ <= $random;
		injection_channels_10_ <= $random;
		injection_channels_9_ <= $random;
		injection_channels_8_ <= $random;
		injection_channels_7_ <= $random;
		injection_channels_6_ <= $random;
		injection_channels_5_ <= $random;
		injection_channels_4_ <= $random;
		injection_channels_3_ <= $random;
		injection_channels_2_ <= $random;
		injection_channels_1_ <= $random;
		injection_channels_0_ <= $random;
		ejection_flow_ctrl_26_ <= $random;
		ejection_flow_ctrl_25_ <= $random;
		ejection_flow_ctrl_24_ <= $random;
		ejection_flow_ctrl_23_ <= $random;
		ejection_flow_ctrl_22_ <= $random;
		ejection_flow_ctrl_21_ <= $random;
		ejection_flow_ctrl_20_ <= $random;
		ejection_flow_ctrl_19_ <= $random;
		ejection_flow_ctrl_18_ <= $random;
		ejection_flow_ctrl_17_ <= $random;
		ejection_flow_ctrl_16_ <= $random;
		ejection_flow_ctrl_15_ <= $random;
		ejection_flow_ctrl_14_ <= $random;
		ejection_flow_ctrl_13_ <= $random;
		ejection_flow_ctrl_12_ <= $random;
		ejection_flow_ctrl_11_ <= $random;
		ejection_flow_ctrl_10_ <= $random;
		ejection_flow_ctrl_9_ <= $random;
		ejection_flow_ctrl_8_ <= $random;
		ejection_flow_ctrl_7_ <= $random;
		ejection_flow_ctrl_6_ <= $random;
		ejection_flow_ctrl_5_ <= $random;
		ejection_flow_ctrl_4_ <= $random;
		ejection_flow_ctrl_3_ <= $random;
		ejection_flow_ctrl_2_ <= $random;
		ejection_flow_ctrl_1_ <= $random;
		ejection_flow_ctrl_0_ <= $random;
	end

// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge clk[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else 
begin
			if(!(injection_flow_ctrl_26__gfpga === injection_flow_ctrl_26__bench) && !(injection_flow_ctrl_26__bench === 1'bx)) begin
				injection_flow_ctrl_26__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_26__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_25__gfpga === injection_flow_ctrl_25__bench) && !(injection_flow_ctrl_25__bench === 1'bx)) begin
				injection_flow_ctrl_25__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_25__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_24__gfpga === injection_flow_ctrl_24__bench) && !(injection_flow_ctrl_24__bench === 1'bx)) begin
				injection_flow_ctrl_24__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_24__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_23__gfpga === injection_flow_ctrl_23__bench) && !(injection_flow_ctrl_23__bench === 1'bx)) begin
				injection_flow_ctrl_23__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_23__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_22__gfpga === injection_flow_ctrl_22__bench) && !(injection_flow_ctrl_22__bench === 1'bx)) begin
				injection_flow_ctrl_22__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_22__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_21__gfpga === injection_flow_ctrl_21__bench) && !(injection_flow_ctrl_21__bench === 1'bx)) begin
				injection_flow_ctrl_21__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_21__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_20__gfpga === injection_flow_ctrl_20__bench) && !(injection_flow_ctrl_20__bench === 1'bx)) begin
				injection_flow_ctrl_20__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_20__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_19__gfpga === injection_flow_ctrl_19__bench) && !(injection_flow_ctrl_19__bench === 1'bx)) begin
				injection_flow_ctrl_19__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_19__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_18__gfpga === injection_flow_ctrl_18__bench) && !(injection_flow_ctrl_18__bench === 1'bx)) begin
				injection_flow_ctrl_18__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_18__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_17__gfpga === injection_flow_ctrl_17__bench) && !(injection_flow_ctrl_17__bench === 1'bx)) begin
				injection_flow_ctrl_17__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_17__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_16__gfpga === injection_flow_ctrl_16__bench) && !(injection_flow_ctrl_16__bench === 1'bx)) begin
				injection_flow_ctrl_16__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_16__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_15__gfpga === injection_flow_ctrl_15__bench) && !(injection_flow_ctrl_15__bench === 1'bx)) begin
				injection_flow_ctrl_15__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_15__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_14__gfpga === injection_flow_ctrl_14__bench) && !(injection_flow_ctrl_14__bench === 1'bx)) begin
				injection_flow_ctrl_14__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_14__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_13__gfpga === injection_flow_ctrl_13__bench) && !(injection_flow_ctrl_13__bench === 1'bx)) begin
				injection_flow_ctrl_13__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_13__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_12__gfpga === injection_flow_ctrl_12__bench) && !(injection_flow_ctrl_12__bench === 1'bx)) begin
				injection_flow_ctrl_12__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_12__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_11__gfpga === injection_flow_ctrl_11__bench) && !(injection_flow_ctrl_11__bench === 1'bx)) begin
				injection_flow_ctrl_11__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_11__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_10__gfpga === injection_flow_ctrl_10__bench) && !(injection_flow_ctrl_10__bench === 1'bx)) begin
				injection_flow_ctrl_10__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_10__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_9__gfpga === injection_flow_ctrl_9__bench) && !(injection_flow_ctrl_9__bench === 1'bx)) begin
				injection_flow_ctrl_9__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_9__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_8__gfpga === injection_flow_ctrl_8__bench) && !(injection_flow_ctrl_8__bench === 1'bx)) begin
				injection_flow_ctrl_8__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_8__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_7__gfpga === injection_flow_ctrl_7__bench) && !(injection_flow_ctrl_7__bench === 1'bx)) begin
				injection_flow_ctrl_7__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_7__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_6__gfpga === injection_flow_ctrl_6__bench) && !(injection_flow_ctrl_6__bench === 1'bx)) begin
				injection_flow_ctrl_6__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_6__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_5__gfpga === injection_flow_ctrl_5__bench) && !(injection_flow_ctrl_5__bench === 1'bx)) begin
				injection_flow_ctrl_5__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_5__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_4__gfpga === injection_flow_ctrl_4__bench) && !(injection_flow_ctrl_4__bench === 1'bx)) begin
				injection_flow_ctrl_4__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_4__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_3__gfpga === injection_flow_ctrl_3__bench) && !(injection_flow_ctrl_3__bench === 1'bx)) begin
				injection_flow_ctrl_3__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_3__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_2__gfpga === injection_flow_ctrl_2__bench) && !(injection_flow_ctrl_2__bench === 1'bx)) begin
				injection_flow_ctrl_2__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_2__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_1__gfpga === injection_flow_ctrl_1__bench) && !(injection_flow_ctrl_1__bench === 1'bx)) begin
				injection_flow_ctrl_1__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_1__flag<= 1'b0;
			end
			if(!(injection_flow_ctrl_0__gfpga === injection_flow_ctrl_0__bench) && !(injection_flow_ctrl_0__bench === 1'bx)) begin
				injection_flow_ctrl_0__flag <= 1'b1;
			end else begin
				injection_flow_ctrl_0__flag<= 1'b0;
			end
			if(!(ejection_channels_629__gfpga === ejection_channels_629__bench) && !(ejection_channels_629__bench === 1'bx)) begin
				ejection_channels_629__flag <= 1'b1;
			end else begin
				ejection_channels_629__flag<= 1'b0;
			end
			if(!(ejection_channels_628__gfpga === ejection_channels_628__bench) && !(ejection_channels_628__bench === 1'bx)) begin
				ejection_channels_628__flag <= 1'b1;
			end else begin
				ejection_channels_628__flag<= 1'b0;
			end
			if(!(ejection_channels_627__gfpga === ejection_channels_627__bench) && !(ejection_channels_627__bench === 1'bx)) begin
				ejection_channels_627__flag <= 1'b1;
			end else begin
				ejection_channels_627__flag<= 1'b0;
			end
			if(!(ejection_channels_626__gfpga === ejection_channels_626__bench) && !(ejection_channels_626__bench === 1'bx)) begin
				ejection_channels_626__flag <= 1'b1;
			end else begin
				ejection_channels_626__flag<= 1'b0;
			end
			if(!(ejection_channels_625__gfpga === ejection_channels_625__bench) && !(ejection_channels_625__bench === 1'bx)) begin
				ejection_channels_625__flag <= 1'b1;
			end else begin
				ejection_channels_625__flag<= 1'b0;
			end
			if(!(ejection_channels_624__gfpga === ejection_channels_624__bench) && !(ejection_channels_624__bench === 1'bx)) begin
				ejection_channels_624__flag <= 1'b1;
			end else begin
				ejection_channels_624__flag<= 1'b0;
			end
			if(!(ejection_channels_623__gfpga === ejection_channels_623__bench) && !(ejection_channels_623__bench === 1'bx)) begin
				ejection_channels_623__flag <= 1'b1;
			end else begin
				ejection_channels_623__flag<= 1'b0;
			end
			if(!(ejection_channels_622__gfpga === ejection_channels_622__bench) && !(ejection_channels_622__bench === 1'bx)) begin
				ejection_channels_622__flag <= 1'b1;
			end else begin
				ejection_channels_622__flag<= 1'b0;
			end
			if(!(ejection_channels_621__gfpga === ejection_channels_621__bench) && !(ejection_channels_621__bench === 1'bx)) begin
				ejection_channels_621__flag <= 1'b1;
			end else begin
				ejection_channels_621__flag<= 1'b0;
			end
			if(!(ejection_channels_620__gfpga === ejection_channels_620__bench) && !(ejection_channels_620__bench === 1'bx)) begin
				ejection_channels_620__flag <= 1'b1;
			end else begin
				ejection_channels_620__flag<= 1'b0;
			end
			if(!(ejection_channels_619__gfpga === ejection_channels_619__bench) && !(ejection_channels_619__bench === 1'bx)) begin
				ejection_channels_619__flag <= 1'b1;
			end else begin
				ejection_channels_619__flag<= 1'b0;
			end
			if(!(ejection_channels_618__gfpga === ejection_channels_618__bench) && !(ejection_channels_618__bench === 1'bx)) begin
				ejection_channels_618__flag <= 1'b1;
			end else begin
				ejection_channels_618__flag<= 1'b0;
			end
			if(!(ejection_channels_617__gfpga === ejection_channels_617__bench) && !(ejection_channels_617__bench === 1'bx)) begin
				ejection_channels_617__flag <= 1'b1;
			end else begin
				ejection_channels_617__flag<= 1'b0;
			end
			if(!(ejection_channels_616__gfpga === ejection_channels_616__bench) && !(ejection_channels_616__bench === 1'bx)) begin
				ejection_channels_616__flag <= 1'b1;
			end else begin
				ejection_channels_616__flag<= 1'b0;
			end
			if(!(ejection_channels_615__gfpga === ejection_channels_615__bench) && !(ejection_channels_615__bench === 1'bx)) begin
				ejection_channels_615__flag <= 1'b1;
			end else begin
				ejection_channels_615__flag<= 1'b0;
			end
			if(!(ejection_channels_614__gfpga === ejection_channels_614__bench) && !(ejection_channels_614__bench === 1'bx)) begin
				ejection_channels_614__flag <= 1'b1;
			end else begin
				ejection_channels_614__flag<= 1'b0;
			end
			if(!(ejection_channels_613__gfpga === ejection_channels_613__bench) && !(ejection_channels_613__bench === 1'bx)) begin
				ejection_channels_613__flag <= 1'b1;
			end else begin
				ejection_channels_613__flag<= 1'b0;
			end
			if(!(ejection_channels_612__gfpga === ejection_channels_612__bench) && !(ejection_channels_612__bench === 1'bx)) begin
				ejection_channels_612__flag <= 1'b1;
			end else begin
				ejection_channels_612__flag<= 1'b0;
			end
			if(!(ejection_channels_611__gfpga === ejection_channels_611__bench) && !(ejection_channels_611__bench === 1'bx)) begin
				ejection_channels_611__flag <= 1'b1;
			end else begin
				ejection_channels_611__flag<= 1'b0;
			end
			if(!(ejection_channels_610__gfpga === ejection_channels_610__bench) && !(ejection_channels_610__bench === 1'bx)) begin
				ejection_channels_610__flag <= 1'b1;
			end else begin
				ejection_channels_610__flag<= 1'b0;
			end
			if(!(ejection_channels_609__gfpga === ejection_channels_609__bench) && !(ejection_channels_609__bench === 1'bx)) begin
				ejection_channels_609__flag <= 1'b1;
			end else begin
				ejection_channels_609__flag<= 1'b0;
			end
			if(!(ejection_channels_608__gfpga === ejection_channels_608__bench) && !(ejection_channels_608__bench === 1'bx)) begin
				ejection_channels_608__flag <= 1'b1;
			end else begin
				ejection_channels_608__flag<= 1'b0;
			end
			if(!(ejection_channels_607__gfpga === ejection_channels_607__bench) && !(ejection_channels_607__bench === 1'bx)) begin
				ejection_channels_607__flag <= 1'b1;
			end else begin
				ejection_channels_607__flag<= 1'b0;
			end
			if(!(ejection_channels_606__gfpga === ejection_channels_606__bench) && !(ejection_channels_606__bench === 1'bx)) begin
				ejection_channels_606__flag <= 1'b1;
			end else begin
				ejection_channels_606__flag<= 1'b0;
			end
			if(!(ejection_channels_605__gfpga === ejection_channels_605__bench) && !(ejection_channels_605__bench === 1'bx)) begin
				ejection_channels_605__flag <= 1'b1;
			end else begin
				ejection_channels_605__flag<= 1'b0;
			end
			if(!(ejection_channels_604__gfpga === ejection_channels_604__bench) && !(ejection_channels_604__bench === 1'bx)) begin
				ejection_channels_604__flag <= 1'b1;
			end else begin
				ejection_channels_604__flag<= 1'b0;
			end
			if(!(ejection_channels_603__gfpga === ejection_channels_603__bench) && !(ejection_channels_603__bench === 1'bx)) begin
				ejection_channels_603__flag <= 1'b1;
			end else begin
				ejection_channels_603__flag<= 1'b0;
			end
			if(!(ejection_channels_602__gfpga === ejection_channels_602__bench) && !(ejection_channels_602__bench === 1'bx)) begin
				ejection_channels_602__flag <= 1'b1;
			end else begin
				ejection_channels_602__flag<= 1'b0;
			end
			if(!(ejection_channels_601__gfpga === ejection_channels_601__bench) && !(ejection_channels_601__bench === 1'bx)) begin
				ejection_channels_601__flag <= 1'b1;
			end else begin
				ejection_channels_601__flag<= 1'b0;
			end
			if(!(ejection_channels_600__gfpga === ejection_channels_600__bench) && !(ejection_channels_600__bench === 1'bx)) begin
				ejection_channels_600__flag <= 1'b1;
			end else begin
				ejection_channels_600__flag<= 1'b0;
			end
			if(!(ejection_channels_599__gfpga === ejection_channels_599__bench) && !(ejection_channels_599__bench === 1'bx)) begin
				ejection_channels_599__flag <= 1'b1;
			end else begin
				ejection_channels_599__flag<= 1'b0;
			end
			if(!(ejection_channels_598__gfpga === ejection_channels_598__bench) && !(ejection_channels_598__bench === 1'bx)) begin
				ejection_channels_598__flag <= 1'b1;
			end else begin
				ejection_channels_598__flag<= 1'b0;
			end
			if(!(ejection_channels_597__gfpga === ejection_channels_597__bench) && !(ejection_channels_597__bench === 1'bx)) begin
				ejection_channels_597__flag <= 1'b1;
			end else begin
				ejection_channels_597__flag<= 1'b0;
			end
			if(!(ejection_channels_596__gfpga === ejection_channels_596__bench) && !(ejection_channels_596__bench === 1'bx)) begin
				ejection_channels_596__flag <= 1'b1;
			end else begin
				ejection_channels_596__flag<= 1'b0;
			end
			if(!(ejection_channels_595__gfpga === ejection_channels_595__bench) && !(ejection_channels_595__bench === 1'bx)) begin
				ejection_channels_595__flag <= 1'b1;
			end else begin
				ejection_channels_595__flag<= 1'b0;
			end
			if(!(ejection_channels_594__gfpga === ejection_channels_594__bench) && !(ejection_channels_594__bench === 1'bx)) begin
				ejection_channels_594__flag <= 1'b1;
			end else begin
				ejection_channels_594__flag<= 1'b0;
			end
			if(!(ejection_channels_593__gfpga === ejection_channels_593__bench) && !(ejection_channels_593__bench === 1'bx)) begin
				ejection_channels_593__flag <= 1'b1;
			end else begin
				ejection_channels_593__flag<= 1'b0;
			end
			if(!(ejection_channels_592__gfpga === ejection_channels_592__bench) && !(ejection_channels_592__bench === 1'bx)) begin
				ejection_channels_592__flag <= 1'b1;
			end else begin
				ejection_channels_592__flag<= 1'b0;
			end
			if(!(ejection_channels_591__gfpga === ejection_channels_591__bench) && !(ejection_channels_591__bench === 1'bx)) begin
				ejection_channels_591__flag <= 1'b1;
			end else begin
				ejection_channels_591__flag<= 1'b0;
			end
			if(!(ejection_channels_590__gfpga === ejection_channels_590__bench) && !(ejection_channels_590__bench === 1'bx)) begin
				ejection_channels_590__flag <= 1'b1;
			end else begin
				ejection_channels_590__flag<= 1'b0;
			end
			if(!(ejection_channels_589__gfpga === ejection_channels_589__bench) && !(ejection_channels_589__bench === 1'bx)) begin
				ejection_channels_589__flag <= 1'b1;
			end else begin
				ejection_channels_589__flag<= 1'b0;
			end
			if(!(ejection_channels_588__gfpga === ejection_channels_588__bench) && !(ejection_channels_588__bench === 1'bx)) begin
				ejection_channels_588__flag <= 1'b1;
			end else begin
				ejection_channels_588__flag<= 1'b0;
			end
			if(!(ejection_channels_587__gfpga === ejection_channels_587__bench) && !(ejection_channels_587__bench === 1'bx)) begin
				ejection_channels_587__flag <= 1'b1;
			end else begin
				ejection_channels_587__flag<= 1'b0;
			end
			if(!(ejection_channels_586__gfpga === ejection_channels_586__bench) && !(ejection_channels_586__bench === 1'bx)) begin
				ejection_channels_586__flag <= 1'b1;
			end else begin
				ejection_channels_586__flag<= 1'b0;
			end
			if(!(ejection_channels_585__gfpga === ejection_channels_585__bench) && !(ejection_channels_585__bench === 1'bx)) begin
				ejection_channels_585__flag <= 1'b1;
			end else begin
				ejection_channels_585__flag<= 1'b0;
			end
			if(!(ejection_channels_584__gfpga === ejection_channels_584__bench) && !(ejection_channels_584__bench === 1'bx)) begin
				ejection_channels_584__flag <= 1'b1;
			end else begin
				ejection_channels_584__flag<= 1'b0;
			end
			if(!(ejection_channels_583__gfpga === ejection_channels_583__bench) && !(ejection_channels_583__bench === 1'bx)) begin
				ejection_channels_583__flag <= 1'b1;
			end else begin
				ejection_channels_583__flag<= 1'b0;
			end
			if(!(ejection_channels_582__gfpga === ejection_channels_582__bench) && !(ejection_channels_582__bench === 1'bx)) begin
				ejection_channels_582__flag <= 1'b1;
			end else begin
				ejection_channels_582__flag<= 1'b0;
			end
			if(!(ejection_channels_581__gfpga === ejection_channels_581__bench) && !(ejection_channels_581__bench === 1'bx)) begin
				ejection_channels_581__flag <= 1'b1;
			end else begin
				ejection_channels_581__flag<= 1'b0;
			end
			if(!(ejection_channels_580__gfpga === ejection_channels_580__bench) && !(ejection_channels_580__bench === 1'bx)) begin
				ejection_channels_580__flag <= 1'b1;
			end else begin
				ejection_channels_580__flag<= 1'b0;
			end
			if(!(ejection_channels_579__gfpga === ejection_channels_579__bench) && !(ejection_channels_579__bench === 1'bx)) begin
				ejection_channels_579__flag <= 1'b1;
			end else begin
				ejection_channels_579__flag<= 1'b0;
			end
			if(!(ejection_channels_578__gfpga === ejection_channels_578__bench) && !(ejection_channels_578__bench === 1'bx)) begin
				ejection_channels_578__flag <= 1'b1;
			end else begin
				ejection_channels_578__flag<= 1'b0;
			end
			if(!(ejection_channels_577__gfpga === ejection_channels_577__bench) && !(ejection_channels_577__bench === 1'bx)) begin
				ejection_channels_577__flag <= 1'b1;
			end else begin
				ejection_channels_577__flag<= 1'b0;
			end
			if(!(ejection_channels_576__gfpga === ejection_channels_576__bench) && !(ejection_channels_576__bench === 1'bx)) begin
				ejection_channels_576__flag <= 1'b1;
			end else begin
				ejection_channels_576__flag<= 1'b0;
			end
			if(!(ejection_channels_575__gfpga === ejection_channels_575__bench) && !(ejection_channels_575__bench === 1'bx)) begin
				ejection_channels_575__flag <= 1'b1;
			end else begin
				ejection_channels_575__flag<= 1'b0;
			end
			if(!(ejection_channels_574__gfpga === ejection_channels_574__bench) && !(ejection_channels_574__bench === 1'bx)) begin
				ejection_channels_574__flag <= 1'b1;
			end else begin
				ejection_channels_574__flag<= 1'b0;
			end
			if(!(ejection_channels_573__gfpga === ejection_channels_573__bench) && !(ejection_channels_573__bench === 1'bx)) begin
				ejection_channels_573__flag <= 1'b1;
			end else begin
				ejection_channels_573__flag<= 1'b0;
			end
			if(!(ejection_channels_572__gfpga === ejection_channels_572__bench) && !(ejection_channels_572__bench === 1'bx)) begin
				ejection_channels_572__flag <= 1'b1;
			end else begin
				ejection_channels_572__flag<= 1'b0;
			end
			if(!(ejection_channels_571__gfpga === ejection_channels_571__bench) && !(ejection_channels_571__bench === 1'bx)) begin
				ejection_channels_571__flag <= 1'b1;
			end else begin
				ejection_channels_571__flag<= 1'b0;
			end
			if(!(ejection_channels_570__gfpga === ejection_channels_570__bench) && !(ejection_channels_570__bench === 1'bx)) begin
				ejection_channels_570__flag <= 1'b1;
			end else begin
				ejection_channels_570__flag<= 1'b0;
			end
			if(!(ejection_channels_569__gfpga === ejection_channels_569__bench) && !(ejection_channels_569__bench === 1'bx)) begin
				ejection_channels_569__flag <= 1'b1;
			end else begin
				ejection_channels_569__flag<= 1'b0;
			end
			if(!(ejection_channels_568__gfpga === ejection_channels_568__bench) && !(ejection_channels_568__bench === 1'bx)) begin
				ejection_channels_568__flag <= 1'b1;
			end else begin
				ejection_channels_568__flag<= 1'b0;
			end
			if(!(ejection_channels_567__gfpga === ejection_channels_567__bench) && !(ejection_channels_567__bench === 1'bx)) begin
				ejection_channels_567__flag <= 1'b1;
			end else begin
				ejection_channels_567__flag<= 1'b0;
			end
			if(!(ejection_channels_566__gfpga === ejection_channels_566__bench) && !(ejection_channels_566__bench === 1'bx)) begin
				ejection_channels_566__flag <= 1'b1;
			end else begin
				ejection_channels_566__flag<= 1'b0;
			end
			if(!(ejection_channels_565__gfpga === ejection_channels_565__bench) && !(ejection_channels_565__bench === 1'bx)) begin
				ejection_channels_565__flag <= 1'b1;
			end else begin
				ejection_channels_565__flag<= 1'b0;
			end
			if(!(ejection_channels_564__gfpga === ejection_channels_564__bench) && !(ejection_channels_564__bench === 1'bx)) begin
				ejection_channels_564__flag <= 1'b1;
			end else begin
				ejection_channels_564__flag<= 1'b0;
			end
			if(!(ejection_channels_563__gfpga === ejection_channels_563__bench) && !(ejection_channels_563__bench === 1'bx)) begin
				ejection_channels_563__flag <= 1'b1;
			end else begin
				ejection_channels_563__flag<= 1'b0;
			end
			if(!(ejection_channels_562__gfpga === ejection_channels_562__bench) && !(ejection_channels_562__bench === 1'bx)) begin
				ejection_channels_562__flag <= 1'b1;
			end else begin
				ejection_channels_562__flag<= 1'b0;
			end
			if(!(ejection_channels_561__gfpga === ejection_channels_561__bench) && !(ejection_channels_561__bench === 1'bx)) begin
				ejection_channels_561__flag <= 1'b1;
			end else begin
				ejection_channels_561__flag<= 1'b0;
			end
			if(!(ejection_channels_560__gfpga === ejection_channels_560__bench) && !(ejection_channels_560__bench === 1'bx)) begin
				ejection_channels_560__flag <= 1'b1;
			end else begin
				ejection_channels_560__flag<= 1'b0;
			end
			if(!(ejection_channels_559__gfpga === ejection_channels_559__bench) && !(ejection_channels_559__bench === 1'bx)) begin
				ejection_channels_559__flag <= 1'b1;
			end else begin
				ejection_channels_559__flag<= 1'b0;
			end
			if(!(ejection_channels_558__gfpga === ejection_channels_558__bench) && !(ejection_channels_558__bench === 1'bx)) begin
				ejection_channels_558__flag <= 1'b1;
			end else begin
				ejection_channels_558__flag<= 1'b0;
			end
			if(!(ejection_channels_557__gfpga === ejection_channels_557__bench) && !(ejection_channels_557__bench === 1'bx)) begin
				ejection_channels_557__flag <= 1'b1;
			end else begin
				ejection_channels_557__flag<= 1'b0;
			end
			if(!(ejection_channels_556__gfpga === ejection_channels_556__bench) && !(ejection_channels_556__bench === 1'bx)) begin
				ejection_channels_556__flag <= 1'b1;
			end else begin
				ejection_channels_556__flag<= 1'b0;
			end
			if(!(ejection_channels_555__gfpga === ejection_channels_555__bench) && !(ejection_channels_555__bench === 1'bx)) begin
				ejection_channels_555__flag <= 1'b1;
			end else begin
				ejection_channels_555__flag<= 1'b0;
			end
			if(!(ejection_channels_554__gfpga === ejection_channels_554__bench) && !(ejection_channels_554__bench === 1'bx)) begin
				ejection_channels_554__flag <= 1'b1;
			end else begin
				ejection_channels_554__flag<= 1'b0;
			end
			if(!(ejection_channels_553__gfpga === ejection_channels_553__bench) && !(ejection_channels_553__bench === 1'bx)) begin
				ejection_channels_553__flag <= 1'b1;
			end else begin
				ejection_channels_553__flag<= 1'b0;
			end
			if(!(ejection_channels_552__gfpga === ejection_channels_552__bench) && !(ejection_channels_552__bench === 1'bx)) begin
				ejection_channels_552__flag <= 1'b1;
			end else begin
				ejection_channels_552__flag<= 1'b0;
			end
			if(!(ejection_channels_551__gfpga === ejection_channels_551__bench) && !(ejection_channels_551__bench === 1'bx)) begin
				ejection_channels_551__flag <= 1'b1;
			end else begin
				ejection_channels_551__flag<= 1'b0;
			end
			if(!(ejection_channels_550__gfpga === ejection_channels_550__bench) && !(ejection_channels_550__bench === 1'bx)) begin
				ejection_channels_550__flag <= 1'b1;
			end else begin
				ejection_channels_550__flag<= 1'b0;
			end
			if(!(ejection_channels_549__gfpga === ejection_channels_549__bench) && !(ejection_channels_549__bench === 1'bx)) begin
				ejection_channels_549__flag <= 1'b1;
			end else begin
				ejection_channels_549__flag<= 1'b0;
			end
			if(!(ejection_channels_548__gfpga === ejection_channels_548__bench) && !(ejection_channels_548__bench === 1'bx)) begin
				ejection_channels_548__flag <= 1'b1;
			end else begin
				ejection_channels_548__flag<= 1'b0;
			end
			if(!(ejection_channels_547__gfpga === ejection_channels_547__bench) && !(ejection_channels_547__bench === 1'bx)) begin
				ejection_channels_547__flag <= 1'b1;
			end else begin
				ejection_channels_547__flag<= 1'b0;
			end
			if(!(ejection_channels_546__gfpga === ejection_channels_546__bench) && !(ejection_channels_546__bench === 1'bx)) begin
				ejection_channels_546__flag <= 1'b1;
			end else begin
				ejection_channels_546__flag<= 1'b0;
			end
			if(!(ejection_channels_545__gfpga === ejection_channels_545__bench) && !(ejection_channels_545__bench === 1'bx)) begin
				ejection_channels_545__flag <= 1'b1;
			end else begin
				ejection_channels_545__flag<= 1'b0;
			end
			if(!(ejection_channels_544__gfpga === ejection_channels_544__bench) && !(ejection_channels_544__bench === 1'bx)) begin
				ejection_channels_544__flag <= 1'b1;
			end else begin
				ejection_channels_544__flag<= 1'b0;
			end
			if(!(ejection_channels_543__gfpga === ejection_channels_543__bench) && !(ejection_channels_543__bench === 1'bx)) begin
				ejection_channels_543__flag <= 1'b1;
			end else begin
				ejection_channels_543__flag<= 1'b0;
			end
			if(!(ejection_channels_542__gfpga === ejection_channels_542__bench) && !(ejection_channels_542__bench === 1'bx)) begin
				ejection_channels_542__flag <= 1'b1;
			end else begin
				ejection_channels_542__flag<= 1'b0;
			end
			if(!(ejection_channels_541__gfpga === ejection_channels_541__bench) && !(ejection_channels_541__bench === 1'bx)) begin
				ejection_channels_541__flag <= 1'b1;
			end else begin
				ejection_channels_541__flag<= 1'b0;
			end
			if(!(ejection_channels_540__gfpga === ejection_channels_540__bench) && !(ejection_channels_540__bench === 1'bx)) begin
				ejection_channels_540__flag <= 1'b1;
			end else begin
				ejection_channels_540__flag<= 1'b0;
			end
			if(!(ejection_channels_539__gfpga === ejection_channels_539__bench) && !(ejection_channels_539__bench === 1'bx)) begin
				ejection_channels_539__flag <= 1'b1;
			end else begin
				ejection_channels_539__flag<= 1'b0;
			end
			if(!(ejection_channels_538__gfpga === ejection_channels_538__bench) && !(ejection_channels_538__bench === 1'bx)) begin
				ejection_channels_538__flag <= 1'b1;
			end else begin
				ejection_channels_538__flag<= 1'b0;
			end
			if(!(ejection_channels_537__gfpga === ejection_channels_537__bench) && !(ejection_channels_537__bench === 1'bx)) begin
				ejection_channels_537__flag <= 1'b1;
			end else begin
				ejection_channels_537__flag<= 1'b0;
			end
			if(!(ejection_channels_536__gfpga === ejection_channels_536__bench) && !(ejection_channels_536__bench === 1'bx)) begin
				ejection_channels_536__flag <= 1'b1;
			end else begin
				ejection_channels_536__flag<= 1'b0;
			end
			if(!(ejection_channels_535__gfpga === ejection_channels_535__bench) && !(ejection_channels_535__bench === 1'bx)) begin
				ejection_channels_535__flag <= 1'b1;
			end else begin
				ejection_channels_535__flag<= 1'b0;
			end
			if(!(ejection_channels_534__gfpga === ejection_channels_534__bench) && !(ejection_channels_534__bench === 1'bx)) begin
				ejection_channels_534__flag <= 1'b1;
			end else begin
				ejection_channels_534__flag<= 1'b0;
			end
			if(!(ejection_channels_533__gfpga === ejection_channels_533__bench) && !(ejection_channels_533__bench === 1'bx)) begin
				ejection_channels_533__flag <= 1'b1;
			end else begin
				ejection_channels_533__flag<= 1'b0;
			end
			if(!(ejection_channels_532__gfpga === ejection_channels_532__bench) && !(ejection_channels_532__bench === 1'bx)) begin
				ejection_channels_532__flag <= 1'b1;
			end else begin
				ejection_channels_532__flag<= 1'b0;
			end
			if(!(ejection_channels_531__gfpga === ejection_channels_531__bench) && !(ejection_channels_531__bench === 1'bx)) begin
				ejection_channels_531__flag <= 1'b1;
			end else begin
				ejection_channels_531__flag<= 1'b0;
			end
			if(!(ejection_channels_530__gfpga === ejection_channels_530__bench) && !(ejection_channels_530__bench === 1'bx)) begin
				ejection_channels_530__flag <= 1'b1;
			end else begin
				ejection_channels_530__flag<= 1'b0;
			end
			if(!(ejection_channels_529__gfpga === ejection_channels_529__bench) && !(ejection_channels_529__bench === 1'bx)) begin
				ejection_channels_529__flag <= 1'b1;
			end else begin
				ejection_channels_529__flag<= 1'b0;
			end
			if(!(ejection_channels_528__gfpga === ejection_channels_528__bench) && !(ejection_channels_528__bench === 1'bx)) begin
				ejection_channels_528__flag <= 1'b1;
			end else begin
				ejection_channels_528__flag<= 1'b0;
			end
			if(!(ejection_channels_527__gfpga === ejection_channels_527__bench) && !(ejection_channels_527__bench === 1'bx)) begin
				ejection_channels_527__flag <= 1'b1;
			end else begin
				ejection_channels_527__flag<= 1'b0;
			end
			if(!(ejection_channels_526__gfpga === ejection_channels_526__bench) && !(ejection_channels_526__bench === 1'bx)) begin
				ejection_channels_526__flag <= 1'b1;
			end else begin
				ejection_channels_526__flag<= 1'b0;
			end
			if(!(ejection_channels_525__gfpga === ejection_channels_525__bench) && !(ejection_channels_525__bench === 1'bx)) begin
				ejection_channels_525__flag <= 1'b1;
			end else begin
				ejection_channels_525__flag<= 1'b0;
			end
			if(!(ejection_channels_524__gfpga === ejection_channels_524__bench) && !(ejection_channels_524__bench === 1'bx)) begin
				ejection_channels_524__flag <= 1'b1;
			end else begin
				ejection_channels_524__flag<= 1'b0;
			end
			if(!(ejection_channels_523__gfpga === ejection_channels_523__bench) && !(ejection_channels_523__bench === 1'bx)) begin
				ejection_channels_523__flag <= 1'b1;
			end else begin
				ejection_channels_523__flag<= 1'b0;
			end
			if(!(ejection_channels_522__gfpga === ejection_channels_522__bench) && !(ejection_channels_522__bench === 1'bx)) begin
				ejection_channels_522__flag <= 1'b1;
			end else begin
				ejection_channels_522__flag<= 1'b0;
			end
			if(!(ejection_channels_521__gfpga === ejection_channels_521__bench) && !(ejection_channels_521__bench === 1'bx)) begin
				ejection_channels_521__flag <= 1'b1;
			end else begin
				ejection_channels_521__flag<= 1'b0;
			end
			if(!(ejection_channels_520__gfpga === ejection_channels_520__bench) && !(ejection_channels_520__bench === 1'bx)) begin
				ejection_channels_520__flag <= 1'b1;
			end else begin
				ejection_channels_520__flag<= 1'b0;
			end
			if(!(ejection_channels_519__gfpga === ejection_channels_519__bench) && !(ejection_channels_519__bench === 1'bx)) begin
				ejection_channels_519__flag <= 1'b1;
			end else begin
				ejection_channels_519__flag<= 1'b0;
			end
			if(!(ejection_channels_518__gfpga === ejection_channels_518__bench) && !(ejection_channels_518__bench === 1'bx)) begin
				ejection_channels_518__flag <= 1'b1;
			end else begin
				ejection_channels_518__flag<= 1'b0;
			end
			if(!(ejection_channels_517__gfpga === ejection_channels_517__bench) && !(ejection_channels_517__bench === 1'bx)) begin
				ejection_channels_517__flag <= 1'b1;
			end else begin
				ejection_channels_517__flag<= 1'b0;
			end
			if(!(ejection_channels_516__gfpga === ejection_channels_516__bench) && !(ejection_channels_516__bench === 1'bx)) begin
				ejection_channels_516__flag <= 1'b1;
			end else begin
				ejection_channels_516__flag<= 1'b0;
			end
			if(!(ejection_channels_515__gfpga === ejection_channels_515__bench) && !(ejection_channels_515__bench === 1'bx)) begin
				ejection_channels_515__flag <= 1'b1;
			end else begin
				ejection_channels_515__flag<= 1'b0;
			end
			if(!(ejection_channels_514__gfpga === ejection_channels_514__bench) && !(ejection_channels_514__bench === 1'bx)) begin
				ejection_channels_514__flag <= 1'b1;
			end else begin
				ejection_channels_514__flag<= 1'b0;
			end
			if(!(ejection_channels_513__gfpga === ejection_channels_513__bench) && !(ejection_channels_513__bench === 1'bx)) begin
				ejection_channels_513__flag <= 1'b1;
			end else begin
				ejection_channels_513__flag<= 1'b0;
			end
			if(!(ejection_channels_512__gfpga === ejection_channels_512__bench) && !(ejection_channels_512__bench === 1'bx)) begin
				ejection_channels_512__flag <= 1'b1;
			end else begin
				ejection_channels_512__flag<= 1'b0;
			end
			if(!(ejection_channels_511__gfpga === ejection_channels_511__bench) && !(ejection_channels_511__bench === 1'bx)) begin
				ejection_channels_511__flag <= 1'b1;
			end else begin
				ejection_channels_511__flag<= 1'b0;
			end
			if(!(ejection_channels_510__gfpga === ejection_channels_510__bench) && !(ejection_channels_510__bench === 1'bx)) begin
				ejection_channels_510__flag <= 1'b1;
			end else begin
				ejection_channels_510__flag<= 1'b0;
			end
			if(!(ejection_channels_509__gfpga === ejection_channels_509__bench) && !(ejection_channels_509__bench === 1'bx)) begin
				ejection_channels_509__flag <= 1'b1;
			end else begin
				ejection_channels_509__flag<= 1'b0;
			end
			if(!(ejection_channels_508__gfpga === ejection_channels_508__bench) && !(ejection_channels_508__bench === 1'bx)) begin
				ejection_channels_508__flag <= 1'b1;
			end else begin
				ejection_channels_508__flag<= 1'b0;
			end
			if(!(ejection_channels_507__gfpga === ejection_channels_507__bench) && !(ejection_channels_507__bench === 1'bx)) begin
				ejection_channels_507__flag <= 1'b1;
			end else begin
				ejection_channels_507__flag<= 1'b0;
			end
			if(!(ejection_channels_506__gfpga === ejection_channels_506__bench) && !(ejection_channels_506__bench === 1'bx)) begin
				ejection_channels_506__flag <= 1'b1;
			end else begin
				ejection_channels_506__flag<= 1'b0;
			end
			if(!(ejection_channels_505__gfpga === ejection_channels_505__bench) && !(ejection_channels_505__bench === 1'bx)) begin
				ejection_channels_505__flag <= 1'b1;
			end else begin
				ejection_channels_505__flag<= 1'b0;
			end
			if(!(ejection_channels_504__gfpga === ejection_channels_504__bench) && !(ejection_channels_504__bench === 1'bx)) begin
				ejection_channels_504__flag <= 1'b1;
			end else begin
				ejection_channels_504__flag<= 1'b0;
			end
			if(!(ejection_channels_503__gfpga === ejection_channels_503__bench) && !(ejection_channels_503__bench === 1'bx)) begin
				ejection_channels_503__flag <= 1'b1;
			end else begin
				ejection_channels_503__flag<= 1'b0;
			end
			if(!(ejection_channels_502__gfpga === ejection_channels_502__bench) && !(ejection_channels_502__bench === 1'bx)) begin
				ejection_channels_502__flag <= 1'b1;
			end else begin
				ejection_channels_502__flag<= 1'b0;
			end
			if(!(ejection_channels_501__gfpga === ejection_channels_501__bench) && !(ejection_channels_501__bench === 1'bx)) begin
				ejection_channels_501__flag <= 1'b1;
			end else begin
				ejection_channels_501__flag<= 1'b0;
			end
			if(!(ejection_channels_500__gfpga === ejection_channels_500__bench) && !(ejection_channels_500__bench === 1'bx)) begin
				ejection_channels_500__flag <= 1'b1;
			end else begin
				ejection_channels_500__flag<= 1'b0;
			end
			if(!(ejection_channels_499__gfpga === ejection_channels_499__bench) && !(ejection_channels_499__bench === 1'bx)) begin
				ejection_channels_499__flag <= 1'b1;
			end else begin
				ejection_channels_499__flag<= 1'b0;
			end
			if(!(ejection_channels_498__gfpga === ejection_channels_498__bench) && !(ejection_channels_498__bench === 1'bx)) begin
				ejection_channels_498__flag <= 1'b1;
			end else begin
				ejection_channels_498__flag<= 1'b0;
			end
			if(!(ejection_channels_497__gfpga === ejection_channels_497__bench) && !(ejection_channels_497__bench === 1'bx)) begin
				ejection_channels_497__flag <= 1'b1;
			end else begin
				ejection_channels_497__flag<= 1'b0;
			end
			if(!(ejection_channels_496__gfpga === ejection_channels_496__bench) && !(ejection_channels_496__bench === 1'bx)) begin
				ejection_channels_496__flag <= 1'b1;
			end else begin
				ejection_channels_496__flag<= 1'b0;
			end
			if(!(ejection_channels_495__gfpga === ejection_channels_495__bench) && !(ejection_channels_495__bench === 1'bx)) begin
				ejection_channels_495__flag <= 1'b1;
			end else begin
				ejection_channels_495__flag<= 1'b0;
			end
			if(!(ejection_channels_494__gfpga === ejection_channels_494__bench) && !(ejection_channels_494__bench === 1'bx)) begin
				ejection_channels_494__flag <= 1'b1;
			end else begin
				ejection_channels_494__flag<= 1'b0;
			end
			if(!(ejection_channels_493__gfpga === ejection_channels_493__bench) && !(ejection_channels_493__bench === 1'bx)) begin
				ejection_channels_493__flag <= 1'b1;
			end else begin
				ejection_channels_493__flag<= 1'b0;
			end
			if(!(ejection_channels_492__gfpga === ejection_channels_492__bench) && !(ejection_channels_492__bench === 1'bx)) begin
				ejection_channels_492__flag <= 1'b1;
			end else begin
				ejection_channels_492__flag<= 1'b0;
			end
			if(!(ejection_channels_491__gfpga === ejection_channels_491__bench) && !(ejection_channels_491__bench === 1'bx)) begin
				ejection_channels_491__flag <= 1'b1;
			end else begin
				ejection_channels_491__flag<= 1'b0;
			end
			if(!(ejection_channels_490__gfpga === ejection_channels_490__bench) && !(ejection_channels_490__bench === 1'bx)) begin
				ejection_channels_490__flag <= 1'b1;
			end else begin
				ejection_channels_490__flag<= 1'b0;
			end
			if(!(ejection_channels_489__gfpga === ejection_channels_489__bench) && !(ejection_channels_489__bench === 1'bx)) begin
				ejection_channels_489__flag <= 1'b1;
			end else begin
				ejection_channels_489__flag<= 1'b0;
			end
			if(!(ejection_channels_488__gfpga === ejection_channels_488__bench) && !(ejection_channels_488__bench === 1'bx)) begin
				ejection_channels_488__flag <= 1'b1;
			end else begin
				ejection_channels_488__flag<= 1'b0;
			end
			if(!(ejection_channels_487__gfpga === ejection_channels_487__bench) && !(ejection_channels_487__bench === 1'bx)) begin
				ejection_channels_487__flag <= 1'b1;
			end else begin
				ejection_channels_487__flag<= 1'b0;
			end
			if(!(ejection_channels_486__gfpga === ejection_channels_486__bench) && !(ejection_channels_486__bench === 1'bx)) begin
				ejection_channels_486__flag <= 1'b1;
			end else begin
				ejection_channels_486__flag<= 1'b0;
			end
			if(!(ejection_channels_485__gfpga === ejection_channels_485__bench) && !(ejection_channels_485__bench === 1'bx)) begin
				ejection_channels_485__flag <= 1'b1;
			end else begin
				ejection_channels_485__flag<= 1'b0;
			end
			if(!(ejection_channels_484__gfpga === ejection_channels_484__bench) && !(ejection_channels_484__bench === 1'bx)) begin
				ejection_channels_484__flag <= 1'b1;
			end else begin
				ejection_channels_484__flag<= 1'b0;
			end
			if(!(ejection_channels_483__gfpga === ejection_channels_483__bench) && !(ejection_channels_483__bench === 1'bx)) begin
				ejection_channels_483__flag <= 1'b1;
			end else begin
				ejection_channels_483__flag<= 1'b0;
			end
			if(!(ejection_channels_482__gfpga === ejection_channels_482__bench) && !(ejection_channels_482__bench === 1'bx)) begin
				ejection_channels_482__flag <= 1'b1;
			end else begin
				ejection_channels_482__flag<= 1'b0;
			end
			if(!(ejection_channels_481__gfpga === ejection_channels_481__bench) && !(ejection_channels_481__bench === 1'bx)) begin
				ejection_channels_481__flag <= 1'b1;
			end else begin
				ejection_channels_481__flag<= 1'b0;
			end
			if(!(ejection_channels_480__gfpga === ejection_channels_480__bench) && !(ejection_channels_480__bench === 1'bx)) begin
				ejection_channels_480__flag <= 1'b1;
			end else begin
				ejection_channels_480__flag<= 1'b0;
			end
			if(!(ejection_channels_479__gfpga === ejection_channels_479__bench) && !(ejection_channels_479__bench === 1'bx)) begin
				ejection_channels_479__flag <= 1'b1;
			end else begin
				ejection_channels_479__flag<= 1'b0;
			end
			if(!(ejection_channels_478__gfpga === ejection_channels_478__bench) && !(ejection_channels_478__bench === 1'bx)) begin
				ejection_channels_478__flag <= 1'b1;
			end else begin
				ejection_channels_478__flag<= 1'b0;
			end
			if(!(ejection_channels_477__gfpga === ejection_channels_477__bench) && !(ejection_channels_477__bench === 1'bx)) begin
				ejection_channels_477__flag <= 1'b1;
			end else begin
				ejection_channels_477__flag<= 1'b0;
			end
			if(!(ejection_channels_476__gfpga === ejection_channels_476__bench) && !(ejection_channels_476__bench === 1'bx)) begin
				ejection_channels_476__flag <= 1'b1;
			end else begin
				ejection_channels_476__flag<= 1'b0;
			end
			if(!(ejection_channels_475__gfpga === ejection_channels_475__bench) && !(ejection_channels_475__bench === 1'bx)) begin
				ejection_channels_475__flag <= 1'b1;
			end else begin
				ejection_channels_475__flag<= 1'b0;
			end
			if(!(ejection_channels_474__gfpga === ejection_channels_474__bench) && !(ejection_channels_474__bench === 1'bx)) begin
				ejection_channels_474__flag <= 1'b1;
			end else begin
				ejection_channels_474__flag<= 1'b0;
			end
			if(!(ejection_channels_473__gfpga === ejection_channels_473__bench) && !(ejection_channels_473__bench === 1'bx)) begin
				ejection_channels_473__flag <= 1'b1;
			end else begin
				ejection_channels_473__flag<= 1'b0;
			end
			if(!(ejection_channels_472__gfpga === ejection_channels_472__bench) && !(ejection_channels_472__bench === 1'bx)) begin
				ejection_channels_472__flag <= 1'b1;
			end else begin
				ejection_channels_472__flag<= 1'b0;
			end
			if(!(ejection_channels_471__gfpga === ejection_channels_471__bench) && !(ejection_channels_471__bench === 1'bx)) begin
				ejection_channels_471__flag <= 1'b1;
			end else begin
				ejection_channels_471__flag<= 1'b0;
			end
			if(!(ejection_channels_470__gfpga === ejection_channels_470__bench) && !(ejection_channels_470__bench === 1'bx)) begin
				ejection_channels_470__flag <= 1'b1;
			end else begin
				ejection_channels_470__flag<= 1'b0;
			end
			if(!(ejection_channels_469__gfpga === ejection_channels_469__bench) && !(ejection_channels_469__bench === 1'bx)) begin
				ejection_channels_469__flag <= 1'b1;
			end else begin
				ejection_channels_469__flag<= 1'b0;
			end
			if(!(ejection_channels_468__gfpga === ejection_channels_468__bench) && !(ejection_channels_468__bench === 1'bx)) begin
				ejection_channels_468__flag <= 1'b1;
			end else begin
				ejection_channels_468__flag<= 1'b0;
			end
			if(!(ejection_channels_467__gfpga === ejection_channels_467__bench) && !(ejection_channels_467__bench === 1'bx)) begin
				ejection_channels_467__flag <= 1'b1;
			end else begin
				ejection_channels_467__flag<= 1'b0;
			end
			if(!(ejection_channels_466__gfpga === ejection_channels_466__bench) && !(ejection_channels_466__bench === 1'bx)) begin
				ejection_channels_466__flag <= 1'b1;
			end else begin
				ejection_channels_466__flag<= 1'b0;
			end
			if(!(ejection_channels_465__gfpga === ejection_channels_465__bench) && !(ejection_channels_465__bench === 1'bx)) begin
				ejection_channels_465__flag <= 1'b1;
			end else begin
				ejection_channels_465__flag<= 1'b0;
			end
			if(!(ejection_channels_464__gfpga === ejection_channels_464__bench) && !(ejection_channels_464__bench === 1'bx)) begin
				ejection_channels_464__flag <= 1'b1;
			end else begin
				ejection_channels_464__flag<= 1'b0;
			end
			if(!(ejection_channels_463__gfpga === ejection_channels_463__bench) && !(ejection_channels_463__bench === 1'bx)) begin
				ejection_channels_463__flag <= 1'b1;
			end else begin
				ejection_channels_463__flag<= 1'b0;
			end
			if(!(ejection_channels_462__gfpga === ejection_channels_462__bench) && !(ejection_channels_462__bench === 1'bx)) begin
				ejection_channels_462__flag <= 1'b1;
			end else begin
				ejection_channels_462__flag<= 1'b0;
			end
			if(!(ejection_channels_461__gfpga === ejection_channels_461__bench) && !(ejection_channels_461__bench === 1'bx)) begin
				ejection_channels_461__flag <= 1'b1;
			end else begin
				ejection_channels_461__flag<= 1'b0;
			end
			if(!(ejection_channels_460__gfpga === ejection_channels_460__bench) && !(ejection_channels_460__bench === 1'bx)) begin
				ejection_channels_460__flag <= 1'b1;
			end else begin
				ejection_channels_460__flag<= 1'b0;
			end
			if(!(ejection_channels_459__gfpga === ejection_channels_459__bench) && !(ejection_channels_459__bench === 1'bx)) begin
				ejection_channels_459__flag <= 1'b1;
			end else begin
				ejection_channels_459__flag<= 1'b0;
			end
			if(!(ejection_channels_458__gfpga === ejection_channels_458__bench) && !(ejection_channels_458__bench === 1'bx)) begin
				ejection_channels_458__flag <= 1'b1;
			end else begin
				ejection_channels_458__flag<= 1'b0;
			end
			if(!(ejection_channels_457__gfpga === ejection_channels_457__bench) && !(ejection_channels_457__bench === 1'bx)) begin
				ejection_channels_457__flag <= 1'b1;
			end else begin
				ejection_channels_457__flag<= 1'b0;
			end
			if(!(ejection_channels_456__gfpga === ejection_channels_456__bench) && !(ejection_channels_456__bench === 1'bx)) begin
				ejection_channels_456__flag <= 1'b1;
			end else begin
				ejection_channels_456__flag<= 1'b0;
			end
			if(!(ejection_channels_455__gfpga === ejection_channels_455__bench) && !(ejection_channels_455__bench === 1'bx)) begin
				ejection_channels_455__flag <= 1'b1;
			end else begin
				ejection_channels_455__flag<= 1'b0;
			end
			if(!(ejection_channels_454__gfpga === ejection_channels_454__bench) && !(ejection_channels_454__bench === 1'bx)) begin
				ejection_channels_454__flag <= 1'b1;
			end else begin
				ejection_channels_454__flag<= 1'b0;
			end
			if(!(ejection_channels_453__gfpga === ejection_channels_453__bench) && !(ejection_channels_453__bench === 1'bx)) begin
				ejection_channels_453__flag <= 1'b1;
			end else begin
				ejection_channels_453__flag<= 1'b0;
			end
			if(!(ejection_channels_452__gfpga === ejection_channels_452__bench) && !(ejection_channels_452__bench === 1'bx)) begin
				ejection_channels_452__flag <= 1'b1;
			end else begin
				ejection_channels_452__flag<= 1'b0;
			end
			if(!(ejection_channels_451__gfpga === ejection_channels_451__bench) && !(ejection_channels_451__bench === 1'bx)) begin
				ejection_channels_451__flag <= 1'b1;
			end else begin
				ejection_channels_451__flag<= 1'b0;
			end
			if(!(ejection_channels_450__gfpga === ejection_channels_450__bench) && !(ejection_channels_450__bench === 1'bx)) begin
				ejection_channels_450__flag <= 1'b1;
			end else begin
				ejection_channels_450__flag<= 1'b0;
			end
			if(!(ejection_channels_449__gfpga === ejection_channels_449__bench) && !(ejection_channels_449__bench === 1'bx)) begin
				ejection_channels_449__flag <= 1'b1;
			end else begin
				ejection_channels_449__flag<= 1'b0;
			end
			if(!(ejection_channels_448__gfpga === ejection_channels_448__bench) && !(ejection_channels_448__bench === 1'bx)) begin
				ejection_channels_448__flag <= 1'b1;
			end else begin
				ejection_channels_448__flag<= 1'b0;
			end
			if(!(ejection_channels_447__gfpga === ejection_channels_447__bench) && !(ejection_channels_447__bench === 1'bx)) begin
				ejection_channels_447__flag <= 1'b1;
			end else begin
				ejection_channels_447__flag<= 1'b0;
			end
			if(!(ejection_channels_446__gfpga === ejection_channels_446__bench) && !(ejection_channels_446__bench === 1'bx)) begin
				ejection_channels_446__flag <= 1'b1;
			end else begin
				ejection_channels_446__flag<= 1'b0;
			end
			if(!(ejection_channels_445__gfpga === ejection_channels_445__bench) && !(ejection_channels_445__bench === 1'bx)) begin
				ejection_channels_445__flag <= 1'b1;
			end else begin
				ejection_channels_445__flag<= 1'b0;
			end
			if(!(ejection_channels_444__gfpga === ejection_channels_444__bench) && !(ejection_channels_444__bench === 1'bx)) begin
				ejection_channels_444__flag <= 1'b1;
			end else begin
				ejection_channels_444__flag<= 1'b0;
			end
			if(!(ejection_channels_443__gfpga === ejection_channels_443__bench) && !(ejection_channels_443__bench === 1'bx)) begin
				ejection_channels_443__flag <= 1'b1;
			end else begin
				ejection_channels_443__flag<= 1'b0;
			end
			if(!(ejection_channels_442__gfpga === ejection_channels_442__bench) && !(ejection_channels_442__bench === 1'bx)) begin
				ejection_channels_442__flag <= 1'b1;
			end else begin
				ejection_channels_442__flag<= 1'b0;
			end
			if(!(ejection_channels_441__gfpga === ejection_channels_441__bench) && !(ejection_channels_441__bench === 1'bx)) begin
				ejection_channels_441__flag <= 1'b1;
			end else begin
				ejection_channels_441__flag<= 1'b0;
			end
			if(!(ejection_channels_440__gfpga === ejection_channels_440__bench) && !(ejection_channels_440__bench === 1'bx)) begin
				ejection_channels_440__flag <= 1'b1;
			end else begin
				ejection_channels_440__flag<= 1'b0;
			end
			if(!(ejection_channels_439__gfpga === ejection_channels_439__bench) && !(ejection_channels_439__bench === 1'bx)) begin
				ejection_channels_439__flag <= 1'b1;
			end else begin
				ejection_channels_439__flag<= 1'b0;
			end
			if(!(ejection_channels_438__gfpga === ejection_channels_438__bench) && !(ejection_channels_438__bench === 1'bx)) begin
				ejection_channels_438__flag <= 1'b1;
			end else begin
				ejection_channels_438__flag<= 1'b0;
			end
			if(!(ejection_channels_437__gfpga === ejection_channels_437__bench) && !(ejection_channels_437__bench === 1'bx)) begin
				ejection_channels_437__flag <= 1'b1;
			end else begin
				ejection_channels_437__flag<= 1'b0;
			end
			if(!(ejection_channels_436__gfpga === ejection_channels_436__bench) && !(ejection_channels_436__bench === 1'bx)) begin
				ejection_channels_436__flag <= 1'b1;
			end else begin
				ejection_channels_436__flag<= 1'b0;
			end
			if(!(ejection_channels_435__gfpga === ejection_channels_435__bench) && !(ejection_channels_435__bench === 1'bx)) begin
				ejection_channels_435__flag <= 1'b1;
			end else begin
				ejection_channels_435__flag<= 1'b0;
			end
			if(!(ejection_channels_434__gfpga === ejection_channels_434__bench) && !(ejection_channels_434__bench === 1'bx)) begin
				ejection_channels_434__flag <= 1'b1;
			end else begin
				ejection_channels_434__flag<= 1'b0;
			end
			if(!(ejection_channels_433__gfpga === ejection_channels_433__bench) && !(ejection_channels_433__bench === 1'bx)) begin
				ejection_channels_433__flag <= 1'b1;
			end else begin
				ejection_channels_433__flag<= 1'b0;
			end
			if(!(ejection_channels_432__gfpga === ejection_channels_432__bench) && !(ejection_channels_432__bench === 1'bx)) begin
				ejection_channels_432__flag <= 1'b1;
			end else begin
				ejection_channels_432__flag<= 1'b0;
			end
			if(!(ejection_channels_431__gfpga === ejection_channels_431__bench) && !(ejection_channels_431__bench === 1'bx)) begin
				ejection_channels_431__flag <= 1'b1;
			end else begin
				ejection_channels_431__flag<= 1'b0;
			end
			if(!(ejection_channels_430__gfpga === ejection_channels_430__bench) && !(ejection_channels_430__bench === 1'bx)) begin
				ejection_channels_430__flag <= 1'b1;
			end else begin
				ejection_channels_430__flag<= 1'b0;
			end
			if(!(ejection_channels_429__gfpga === ejection_channels_429__bench) && !(ejection_channels_429__bench === 1'bx)) begin
				ejection_channels_429__flag <= 1'b1;
			end else begin
				ejection_channels_429__flag<= 1'b0;
			end
			if(!(ejection_channels_428__gfpga === ejection_channels_428__bench) && !(ejection_channels_428__bench === 1'bx)) begin
				ejection_channels_428__flag <= 1'b1;
			end else begin
				ejection_channels_428__flag<= 1'b0;
			end
			if(!(ejection_channels_427__gfpga === ejection_channels_427__bench) && !(ejection_channels_427__bench === 1'bx)) begin
				ejection_channels_427__flag <= 1'b1;
			end else begin
				ejection_channels_427__flag<= 1'b0;
			end
			if(!(ejection_channels_426__gfpga === ejection_channels_426__bench) && !(ejection_channels_426__bench === 1'bx)) begin
				ejection_channels_426__flag <= 1'b1;
			end else begin
				ejection_channels_426__flag<= 1'b0;
			end
			if(!(ejection_channels_425__gfpga === ejection_channels_425__bench) && !(ejection_channels_425__bench === 1'bx)) begin
				ejection_channels_425__flag <= 1'b1;
			end else begin
				ejection_channels_425__flag<= 1'b0;
			end
			if(!(ejection_channels_424__gfpga === ejection_channels_424__bench) && !(ejection_channels_424__bench === 1'bx)) begin
				ejection_channels_424__flag <= 1'b1;
			end else begin
				ejection_channels_424__flag<= 1'b0;
			end
			if(!(ejection_channels_423__gfpga === ejection_channels_423__bench) && !(ejection_channels_423__bench === 1'bx)) begin
				ejection_channels_423__flag <= 1'b1;
			end else begin
				ejection_channels_423__flag<= 1'b0;
			end
			if(!(ejection_channels_422__gfpga === ejection_channels_422__bench) && !(ejection_channels_422__bench === 1'bx)) begin
				ejection_channels_422__flag <= 1'b1;
			end else begin
				ejection_channels_422__flag<= 1'b0;
			end
			if(!(ejection_channels_421__gfpga === ejection_channels_421__bench) && !(ejection_channels_421__bench === 1'bx)) begin
				ejection_channels_421__flag <= 1'b1;
			end else begin
				ejection_channels_421__flag<= 1'b0;
			end
			if(!(ejection_channels_420__gfpga === ejection_channels_420__bench) && !(ejection_channels_420__bench === 1'bx)) begin
				ejection_channels_420__flag <= 1'b1;
			end else begin
				ejection_channels_420__flag<= 1'b0;
			end
			if(!(ejection_channels_419__gfpga === ejection_channels_419__bench) && !(ejection_channels_419__bench === 1'bx)) begin
				ejection_channels_419__flag <= 1'b1;
			end else begin
				ejection_channels_419__flag<= 1'b0;
			end
			if(!(ejection_channels_418__gfpga === ejection_channels_418__bench) && !(ejection_channels_418__bench === 1'bx)) begin
				ejection_channels_418__flag <= 1'b1;
			end else begin
				ejection_channels_418__flag<= 1'b0;
			end
			if(!(ejection_channels_417__gfpga === ejection_channels_417__bench) && !(ejection_channels_417__bench === 1'bx)) begin
				ejection_channels_417__flag <= 1'b1;
			end else begin
				ejection_channels_417__flag<= 1'b0;
			end
			if(!(ejection_channels_416__gfpga === ejection_channels_416__bench) && !(ejection_channels_416__bench === 1'bx)) begin
				ejection_channels_416__flag <= 1'b1;
			end else begin
				ejection_channels_416__flag<= 1'b0;
			end
			if(!(ejection_channels_415__gfpga === ejection_channels_415__bench) && !(ejection_channels_415__bench === 1'bx)) begin
				ejection_channels_415__flag <= 1'b1;
			end else begin
				ejection_channels_415__flag<= 1'b0;
			end
			if(!(ejection_channels_414__gfpga === ejection_channels_414__bench) && !(ejection_channels_414__bench === 1'bx)) begin
				ejection_channels_414__flag <= 1'b1;
			end else begin
				ejection_channels_414__flag<= 1'b0;
			end
			if(!(ejection_channels_413__gfpga === ejection_channels_413__bench) && !(ejection_channels_413__bench === 1'bx)) begin
				ejection_channels_413__flag <= 1'b1;
			end else begin
				ejection_channels_413__flag<= 1'b0;
			end
			if(!(ejection_channels_412__gfpga === ejection_channels_412__bench) && !(ejection_channels_412__bench === 1'bx)) begin
				ejection_channels_412__flag <= 1'b1;
			end else begin
				ejection_channels_412__flag<= 1'b0;
			end
			if(!(ejection_channels_411__gfpga === ejection_channels_411__bench) && !(ejection_channels_411__bench === 1'bx)) begin
				ejection_channels_411__flag <= 1'b1;
			end else begin
				ejection_channels_411__flag<= 1'b0;
			end
			if(!(ejection_channels_410__gfpga === ejection_channels_410__bench) && !(ejection_channels_410__bench === 1'bx)) begin
				ejection_channels_410__flag <= 1'b1;
			end else begin
				ejection_channels_410__flag<= 1'b0;
			end
			if(!(ejection_channels_409__gfpga === ejection_channels_409__bench) && !(ejection_channels_409__bench === 1'bx)) begin
				ejection_channels_409__flag <= 1'b1;
			end else begin
				ejection_channels_409__flag<= 1'b0;
			end
			if(!(ejection_channels_408__gfpga === ejection_channels_408__bench) && !(ejection_channels_408__bench === 1'bx)) begin
				ejection_channels_408__flag <= 1'b1;
			end else begin
				ejection_channels_408__flag<= 1'b0;
			end
			if(!(ejection_channels_407__gfpga === ejection_channels_407__bench) && !(ejection_channels_407__bench === 1'bx)) begin
				ejection_channels_407__flag <= 1'b1;
			end else begin
				ejection_channels_407__flag<= 1'b0;
			end
			if(!(ejection_channels_406__gfpga === ejection_channels_406__bench) && !(ejection_channels_406__bench === 1'bx)) begin
				ejection_channels_406__flag <= 1'b1;
			end else begin
				ejection_channels_406__flag<= 1'b0;
			end
			if(!(ejection_channels_405__gfpga === ejection_channels_405__bench) && !(ejection_channels_405__bench === 1'bx)) begin
				ejection_channels_405__flag <= 1'b1;
			end else begin
				ejection_channels_405__flag<= 1'b0;
			end
			if(!(ejection_channels_404__gfpga === ejection_channels_404__bench) && !(ejection_channels_404__bench === 1'bx)) begin
				ejection_channels_404__flag <= 1'b1;
			end else begin
				ejection_channels_404__flag<= 1'b0;
			end
			if(!(ejection_channels_403__gfpga === ejection_channels_403__bench) && !(ejection_channels_403__bench === 1'bx)) begin
				ejection_channels_403__flag <= 1'b1;
			end else begin
				ejection_channels_403__flag<= 1'b0;
			end
			if(!(ejection_channels_402__gfpga === ejection_channels_402__bench) && !(ejection_channels_402__bench === 1'bx)) begin
				ejection_channels_402__flag <= 1'b1;
			end else begin
				ejection_channels_402__flag<= 1'b0;
			end
			if(!(ejection_channels_401__gfpga === ejection_channels_401__bench) && !(ejection_channels_401__bench === 1'bx)) begin
				ejection_channels_401__flag <= 1'b1;
			end else begin
				ejection_channels_401__flag<= 1'b0;
			end
			if(!(ejection_channels_400__gfpga === ejection_channels_400__bench) && !(ejection_channels_400__bench === 1'bx)) begin
				ejection_channels_400__flag <= 1'b1;
			end else begin
				ejection_channels_400__flag<= 1'b0;
			end
			if(!(ejection_channels_399__gfpga === ejection_channels_399__bench) && !(ejection_channels_399__bench === 1'bx)) begin
				ejection_channels_399__flag <= 1'b1;
			end else begin
				ejection_channels_399__flag<= 1'b0;
			end
			if(!(ejection_channels_398__gfpga === ejection_channels_398__bench) && !(ejection_channels_398__bench === 1'bx)) begin
				ejection_channels_398__flag <= 1'b1;
			end else begin
				ejection_channels_398__flag<= 1'b0;
			end
			if(!(ejection_channels_397__gfpga === ejection_channels_397__bench) && !(ejection_channels_397__bench === 1'bx)) begin
				ejection_channels_397__flag <= 1'b1;
			end else begin
				ejection_channels_397__flag<= 1'b0;
			end
			if(!(ejection_channels_396__gfpga === ejection_channels_396__bench) && !(ejection_channels_396__bench === 1'bx)) begin
				ejection_channels_396__flag <= 1'b1;
			end else begin
				ejection_channels_396__flag<= 1'b0;
			end
			if(!(ejection_channels_395__gfpga === ejection_channels_395__bench) && !(ejection_channels_395__bench === 1'bx)) begin
				ejection_channels_395__flag <= 1'b1;
			end else begin
				ejection_channels_395__flag<= 1'b0;
			end
			if(!(ejection_channels_394__gfpga === ejection_channels_394__bench) && !(ejection_channels_394__bench === 1'bx)) begin
				ejection_channels_394__flag <= 1'b1;
			end else begin
				ejection_channels_394__flag<= 1'b0;
			end
			if(!(ejection_channels_393__gfpga === ejection_channels_393__bench) && !(ejection_channels_393__bench === 1'bx)) begin
				ejection_channels_393__flag <= 1'b1;
			end else begin
				ejection_channels_393__flag<= 1'b0;
			end
			if(!(ejection_channels_392__gfpga === ejection_channels_392__bench) && !(ejection_channels_392__bench === 1'bx)) begin
				ejection_channels_392__flag <= 1'b1;
			end else begin
				ejection_channels_392__flag<= 1'b0;
			end
			if(!(ejection_channels_391__gfpga === ejection_channels_391__bench) && !(ejection_channels_391__bench === 1'bx)) begin
				ejection_channels_391__flag <= 1'b1;
			end else begin
				ejection_channels_391__flag<= 1'b0;
			end
			if(!(ejection_channels_390__gfpga === ejection_channels_390__bench) && !(ejection_channels_390__bench === 1'bx)) begin
				ejection_channels_390__flag <= 1'b1;
			end else begin
				ejection_channels_390__flag<= 1'b0;
			end
			if(!(ejection_channels_389__gfpga === ejection_channels_389__bench) && !(ejection_channels_389__bench === 1'bx)) begin
				ejection_channels_389__flag <= 1'b1;
			end else begin
				ejection_channels_389__flag<= 1'b0;
			end
			if(!(ejection_channels_388__gfpga === ejection_channels_388__bench) && !(ejection_channels_388__bench === 1'bx)) begin
				ejection_channels_388__flag <= 1'b1;
			end else begin
				ejection_channels_388__flag<= 1'b0;
			end
			if(!(ejection_channels_387__gfpga === ejection_channels_387__bench) && !(ejection_channels_387__bench === 1'bx)) begin
				ejection_channels_387__flag <= 1'b1;
			end else begin
				ejection_channels_387__flag<= 1'b0;
			end
			if(!(ejection_channels_386__gfpga === ejection_channels_386__bench) && !(ejection_channels_386__bench === 1'bx)) begin
				ejection_channels_386__flag <= 1'b1;
			end else begin
				ejection_channels_386__flag<= 1'b0;
			end
			if(!(ejection_channels_385__gfpga === ejection_channels_385__bench) && !(ejection_channels_385__bench === 1'bx)) begin
				ejection_channels_385__flag <= 1'b1;
			end else begin
				ejection_channels_385__flag<= 1'b0;
			end
			if(!(ejection_channels_384__gfpga === ejection_channels_384__bench) && !(ejection_channels_384__bench === 1'bx)) begin
				ejection_channels_384__flag <= 1'b1;
			end else begin
				ejection_channels_384__flag<= 1'b0;
			end
			if(!(ejection_channels_383__gfpga === ejection_channels_383__bench) && !(ejection_channels_383__bench === 1'bx)) begin
				ejection_channels_383__flag <= 1'b1;
			end else begin
				ejection_channels_383__flag<= 1'b0;
			end
			if(!(ejection_channels_382__gfpga === ejection_channels_382__bench) && !(ejection_channels_382__bench === 1'bx)) begin
				ejection_channels_382__flag <= 1'b1;
			end else begin
				ejection_channels_382__flag<= 1'b0;
			end
			if(!(ejection_channels_381__gfpga === ejection_channels_381__bench) && !(ejection_channels_381__bench === 1'bx)) begin
				ejection_channels_381__flag <= 1'b1;
			end else begin
				ejection_channels_381__flag<= 1'b0;
			end
			if(!(ejection_channels_380__gfpga === ejection_channels_380__bench) && !(ejection_channels_380__bench === 1'bx)) begin
				ejection_channels_380__flag <= 1'b1;
			end else begin
				ejection_channels_380__flag<= 1'b0;
			end
			if(!(ejection_channels_379__gfpga === ejection_channels_379__bench) && !(ejection_channels_379__bench === 1'bx)) begin
				ejection_channels_379__flag <= 1'b1;
			end else begin
				ejection_channels_379__flag<= 1'b0;
			end
			if(!(ejection_channels_378__gfpga === ejection_channels_378__bench) && !(ejection_channels_378__bench === 1'bx)) begin
				ejection_channels_378__flag <= 1'b1;
			end else begin
				ejection_channels_378__flag<= 1'b0;
			end
			if(!(ejection_channels_377__gfpga === ejection_channels_377__bench) && !(ejection_channels_377__bench === 1'bx)) begin
				ejection_channels_377__flag <= 1'b1;
			end else begin
				ejection_channels_377__flag<= 1'b0;
			end
			if(!(ejection_channels_376__gfpga === ejection_channels_376__bench) && !(ejection_channels_376__bench === 1'bx)) begin
				ejection_channels_376__flag <= 1'b1;
			end else begin
				ejection_channels_376__flag<= 1'b0;
			end
			if(!(ejection_channels_375__gfpga === ejection_channels_375__bench) && !(ejection_channels_375__bench === 1'bx)) begin
				ejection_channels_375__flag <= 1'b1;
			end else begin
				ejection_channels_375__flag<= 1'b0;
			end
			if(!(ejection_channels_374__gfpga === ejection_channels_374__bench) && !(ejection_channels_374__bench === 1'bx)) begin
				ejection_channels_374__flag <= 1'b1;
			end else begin
				ejection_channels_374__flag<= 1'b0;
			end
			if(!(ejection_channels_373__gfpga === ejection_channels_373__bench) && !(ejection_channels_373__bench === 1'bx)) begin
				ejection_channels_373__flag <= 1'b1;
			end else begin
				ejection_channels_373__flag<= 1'b0;
			end
			if(!(ejection_channels_372__gfpga === ejection_channels_372__bench) && !(ejection_channels_372__bench === 1'bx)) begin
				ejection_channels_372__flag <= 1'b1;
			end else begin
				ejection_channels_372__flag<= 1'b0;
			end
			if(!(ejection_channels_371__gfpga === ejection_channels_371__bench) && !(ejection_channels_371__bench === 1'bx)) begin
				ejection_channels_371__flag <= 1'b1;
			end else begin
				ejection_channels_371__flag<= 1'b0;
			end
			if(!(ejection_channels_370__gfpga === ejection_channels_370__bench) && !(ejection_channels_370__bench === 1'bx)) begin
				ejection_channels_370__flag <= 1'b1;
			end else begin
				ejection_channels_370__flag<= 1'b0;
			end
			if(!(ejection_channels_369__gfpga === ejection_channels_369__bench) && !(ejection_channels_369__bench === 1'bx)) begin
				ejection_channels_369__flag <= 1'b1;
			end else begin
				ejection_channels_369__flag<= 1'b0;
			end
			if(!(ejection_channels_368__gfpga === ejection_channels_368__bench) && !(ejection_channels_368__bench === 1'bx)) begin
				ejection_channels_368__flag <= 1'b1;
			end else begin
				ejection_channels_368__flag<= 1'b0;
			end
			if(!(ejection_channels_367__gfpga === ejection_channels_367__bench) && !(ejection_channels_367__bench === 1'bx)) begin
				ejection_channels_367__flag <= 1'b1;
			end else begin
				ejection_channels_367__flag<= 1'b0;
			end
			if(!(ejection_channels_366__gfpga === ejection_channels_366__bench) && !(ejection_channels_366__bench === 1'bx)) begin
				ejection_channels_366__flag <= 1'b1;
			end else begin
				ejection_channels_366__flag<= 1'b0;
			end
			if(!(ejection_channels_365__gfpga === ejection_channels_365__bench) && !(ejection_channels_365__bench === 1'bx)) begin
				ejection_channels_365__flag <= 1'b1;
			end else begin
				ejection_channels_365__flag<= 1'b0;
			end
			if(!(ejection_channels_364__gfpga === ejection_channels_364__bench) && !(ejection_channels_364__bench === 1'bx)) begin
				ejection_channels_364__flag <= 1'b1;
			end else begin
				ejection_channels_364__flag<= 1'b0;
			end
			if(!(ejection_channels_363__gfpga === ejection_channels_363__bench) && !(ejection_channels_363__bench === 1'bx)) begin
				ejection_channels_363__flag <= 1'b1;
			end else begin
				ejection_channels_363__flag<= 1'b0;
			end
			if(!(ejection_channels_362__gfpga === ejection_channels_362__bench) && !(ejection_channels_362__bench === 1'bx)) begin
				ejection_channels_362__flag <= 1'b1;
			end else begin
				ejection_channels_362__flag<= 1'b0;
			end
			if(!(ejection_channels_361__gfpga === ejection_channels_361__bench) && !(ejection_channels_361__bench === 1'bx)) begin
				ejection_channels_361__flag <= 1'b1;
			end else begin
				ejection_channels_361__flag<= 1'b0;
			end
			if(!(ejection_channels_360__gfpga === ejection_channels_360__bench) && !(ejection_channels_360__bench === 1'bx)) begin
				ejection_channels_360__flag <= 1'b1;
			end else begin
				ejection_channels_360__flag<= 1'b0;
			end
			if(!(ejection_channels_359__gfpga === ejection_channels_359__bench) && !(ejection_channels_359__bench === 1'bx)) begin
				ejection_channels_359__flag <= 1'b1;
			end else begin
				ejection_channels_359__flag<= 1'b0;
			end
			if(!(ejection_channels_358__gfpga === ejection_channels_358__bench) && !(ejection_channels_358__bench === 1'bx)) begin
				ejection_channels_358__flag <= 1'b1;
			end else begin
				ejection_channels_358__flag<= 1'b0;
			end
			if(!(ejection_channels_357__gfpga === ejection_channels_357__bench) && !(ejection_channels_357__bench === 1'bx)) begin
				ejection_channels_357__flag <= 1'b1;
			end else begin
				ejection_channels_357__flag<= 1'b0;
			end
			if(!(ejection_channels_356__gfpga === ejection_channels_356__bench) && !(ejection_channels_356__bench === 1'bx)) begin
				ejection_channels_356__flag <= 1'b1;
			end else begin
				ejection_channels_356__flag<= 1'b0;
			end
			if(!(ejection_channels_355__gfpga === ejection_channels_355__bench) && !(ejection_channels_355__bench === 1'bx)) begin
				ejection_channels_355__flag <= 1'b1;
			end else begin
				ejection_channels_355__flag<= 1'b0;
			end
			if(!(ejection_channels_354__gfpga === ejection_channels_354__bench) && !(ejection_channels_354__bench === 1'bx)) begin
				ejection_channels_354__flag <= 1'b1;
			end else begin
				ejection_channels_354__flag<= 1'b0;
			end
			if(!(ejection_channels_353__gfpga === ejection_channels_353__bench) && !(ejection_channels_353__bench === 1'bx)) begin
				ejection_channels_353__flag <= 1'b1;
			end else begin
				ejection_channels_353__flag<= 1'b0;
			end
			if(!(ejection_channels_352__gfpga === ejection_channels_352__bench) && !(ejection_channels_352__bench === 1'bx)) begin
				ejection_channels_352__flag <= 1'b1;
			end else begin
				ejection_channels_352__flag<= 1'b0;
			end
			if(!(ejection_channels_351__gfpga === ejection_channels_351__bench) && !(ejection_channels_351__bench === 1'bx)) begin
				ejection_channels_351__flag <= 1'b1;
			end else begin
				ejection_channels_351__flag<= 1'b0;
			end
			if(!(ejection_channels_350__gfpga === ejection_channels_350__bench) && !(ejection_channels_350__bench === 1'bx)) begin
				ejection_channels_350__flag <= 1'b1;
			end else begin
				ejection_channels_350__flag<= 1'b0;
			end
			if(!(ejection_channels_349__gfpga === ejection_channels_349__bench) && !(ejection_channels_349__bench === 1'bx)) begin
				ejection_channels_349__flag <= 1'b1;
			end else begin
				ejection_channels_349__flag<= 1'b0;
			end
			if(!(ejection_channels_348__gfpga === ejection_channels_348__bench) && !(ejection_channels_348__bench === 1'bx)) begin
				ejection_channels_348__flag <= 1'b1;
			end else begin
				ejection_channels_348__flag<= 1'b0;
			end
			if(!(ejection_channels_347__gfpga === ejection_channels_347__bench) && !(ejection_channels_347__bench === 1'bx)) begin
				ejection_channels_347__flag <= 1'b1;
			end else begin
				ejection_channels_347__flag<= 1'b0;
			end
			if(!(ejection_channels_346__gfpga === ejection_channels_346__bench) && !(ejection_channels_346__bench === 1'bx)) begin
				ejection_channels_346__flag <= 1'b1;
			end else begin
				ejection_channels_346__flag<= 1'b0;
			end
			if(!(ejection_channels_345__gfpga === ejection_channels_345__bench) && !(ejection_channels_345__bench === 1'bx)) begin
				ejection_channels_345__flag <= 1'b1;
			end else begin
				ejection_channels_345__flag<= 1'b0;
			end
			if(!(ejection_channels_344__gfpga === ejection_channels_344__bench) && !(ejection_channels_344__bench === 1'bx)) begin
				ejection_channels_344__flag <= 1'b1;
			end else begin
				ejection_channels_344__flag<= 1'b0;
			end
			if(!(ejection_channels_343__gfpga === ejection_channels_343__bench) && !(ejection_channels_343__bench === 1'bx)) begin
				ejection_channels_343__flag <= 1'b1;
			end else begin
				ejection_channels_343__flag<= 1'b0;
			end
			if(!(ejection_channels_342__gfpga === ejection_channels_342__bench) && !(ejection_channels_342__bench === 1'bx)) begin
				ejection_channels_342__flag <= 1'b1;
			end else begin
				ejection_channels_342__flag<= 1'b0;
			end
			if(!(ejection_channels_341__gfpga === ejection_channels_341__bench) && !(ejection_channels_341__bench === 1'bx)) begin
				ejection_channels_341__flag <= 1'b1;
			end else begin
				ejection_channels_341__flag<= 1'b0;
			end
			if(!(ejection_channels_340__gfpga === ejection_channels_340__bench) && !(ejection_channels_340__bench === 1'bx)) begin
				ejection_channels_340__flag <= 1'b1;
			end else begin
				ejection_channels_340__flag<= 1'b0;
			end
			if(!(ejection_channels_339__gfpga === ejection_channels_339__bench) && !(ejection_channels_339__bench === 1'bx)) begin
				ejection_channels_339__flag <= 1'b1;
			end else begin
				ejection_channels_339__flag<= 1'b0;
			end
			if(!(ejection_channels_338__gfpga === ejection_channels_338__bench) && !(ejection_channels_338__bench === 1'bx)) begin
				ejection_channels_338__flag <= 1'b1;
			end else begin
				ejection_channels_338__flag<= 1'b0;
			end
			if(!(ejection_channels_337__gfpga === ejection_channels_337__bench) && !(ejection_channels_337__bench === 1'bx)) begin
				ejection_channels_337__flag <= 1'b1;
			end else begin
				ejection_channels_337__flag<= 1'b0;
			end
			if(!(ejection_channels_336__gfpga === ejection_channels_336__bench) && !(ejection_channels_336__bench === 1'bx)) begin
				ejection_channels_336__flag <= 1'b1;
			end else begin
				ejection_channels_336__flag<= 1'b0;
			end
			if(!(ejection_channels_335__gfpga === ejection_channels_335__bench) && !(ejection_channels_335__bench === 1'bx)) begin
				ejection_channels_335__flag <= 1'b1;
			end else begin
				ejection_channels_335__flag<= 1'b0;
			end
			if(!(ejection_channels_334__gfpga === ejection_channels_334__bench) && !(ejection_channels_334__bench === 1'bx)) begin
				ejection_channels_334__flag <= 1'b1;
			end else begin
				ejection_channels_334__flag<= 1'b0;
			end
			if(!(ejection_channels_333__gfpga === ejection_channels_333__bench) && !(ejection_channels_333__bench === 1'bx)) begin
				ejection_channels_333__flag <= 1'b1;
			end else begin
				ejection_channels_333__flag<= 1'b0;
			end
			if(!(ejection_channels_332__gfpga === ejection_channels_332__bench) && !(ejection_channels_332__bench === 1'bx)) begin
				ejection_channels_332__flag <= 1'b1;
			end else begin
				ejection_channels_332__flag<= 1'b0;
			end
			if(!(ejection_channels_331__gfpga === ejection_channels_331__bench) && !(ejection_channels_331__bench === 1'bx)) begin
				ejection_channels_331__flag <= 1'b1;
			end else begin
				ejection_channels_331__flag<= 1'b0;
			end
			if(!(ejection_channels_330__gfpga === ejection_channels_330__bench) && !(ejection_channels_330__bench === 1'bx)) begin
				ejection_channels_330__flag <= 1'b1;
			end else begin
				ejection_channels_330__flag<= 1'b0;
			end
			if(!(ejection_channels_329__gfpga === ejection_channels_329__bench) && !(ejection_channels_329__bench === 1'bx)) begin
				ejection_channels_329__flag <= 1'b1;
			end else begin
				ejection_channels_329__flag<= 1'b0;
			end
			if(!(ejection_channels_328__gfpga === ejection_channels_328__bench) && !(ejection_channels_328__bench === 1'bx)) begin
				ejection_channels_328__flag <= 1'b1;
			end else begin
				ejection_channels_328__flag<= 1'b0;
			end
			if(!(ejection_channels_327__gfpga === ejection_channels_327__bench) && !(ejection_channels_327__bench === 1'bx)) begin
				ejection_channels_327__flag <= 1'b1;
			end else begin
				ejection_channels_327__flag<= 1'b0;
			end
			if(!(ejection_channels_326__gfpga === ejection_channels_326__bench) && !(ejection_channels_326__bench === 1'bx)) begin
				ejection_channels_326__flag <= 1'b1;
			end else begin
				ejection_channels_326__flag<= 1'b0;
			end
			if(!(ejection_channels_325__gfpga === ejection_channels_325__bench) && !(ejection_channels_325__bench === 1'bx)) begin
				ejection_channels_325__flag <= 1'b1;
			end else begin
				ejection_channels_325__flag<= 1'b0;
			end
			if(!(ejection_channels_324__gfpga === ejection_channels_324__bench) && !(ejection_channels_324__bench === 1'bx)) begin
				ejection_channels_324__flag <= 1'b1;
			end else begin
				ejection_channels_324__flag<= 1'b0;
			end
			if(!(ejection_channels_323__gfpga === ejection_channels_323__bench) && !(ejection_channels_323__bench === 1'bx)) begin
				ejection_channels_323__flag <= 1'b1;
			end else begin
				ejection_channels_323__flag<= 1'b0;
			end
			if(!(ejection_channels_322__gfpga === ejection_channels_322__bench) && !(ejection_channels_322__bench === 1'bx)) begin
				ejection_channels_322__flag <= 1'b1;
			end else begin
				ejection_channels_322__flag<= 1'b0;
			end
			if(!(ejection_channels_321__gfpga === ejection_channels_321__bench) && !(ejection_channels_321__bench === 1'bx)) begin
				ejection_channels_321__flag <= 1'b1;
			end else begin
				ejection_channels_321__flag<= 1'b0;
			end
			if(!(ejection_channels_320__gfpga === ejection_channels_320__bench) && !(ejection_channels_320__bench === 1'bx)) begin
				ejection_channels_320__flag <= 1'b1;
			end else begin
				ejection_channels_320__flag<= 1'b0;
			end
			if(!(ejection_channels_319__gfpga === ejection_channels_319__bench) && !(ejection_channels_319__bench === 1'bx)) begin
				ejection_channels_319__flag <= 1'b1;
			end else begin
				ejection_channels_319__flag<= 1'b0;
			end
			if(!(ejection_channels_318__gfpga === ejection_channels_318__bench) && !(ejection_channels_318__bench === 1'bx)) begin
				ejection_channels_318__flag <= 1'b1;
			end else begin
				ejection_channels_318__flag<= 1'b0;
			end
			if(!(ejection_channels_317__gfpga === ejection_channels_317__bench) && !(ejection_channels_317__bench === 1'bx)) begin
				ejection_channels_317__flag <= 1'b1;
			end else begin
				ejection_channels_317__flag<= 1'b0;
			end
			if(!(ejection_channels_316__gfpga === ejection_channels_316__bench) && !(ejection_channels_316__bench === 1'bx)) begin
				ejection_channels_316__flag <= 1'b1;
			end else begin
				ejection_channels_316__flag<= 1'b0;
			end
			if(!(ejection_channels_315__gfpga === ejection_channels_315__bench) && !(ejection_channels_315__bench === 1'bx)) begin
				ejection_channels_315__flag <= 1'b1;
			end else begin
				ejection_channels_315__flag<= 1'b0;
			end
			if(!(ejection_channels_314__gfpga === ejection_channels_314__bench) && !(ejection_channels_314__bench === 1'bx)) begin
				ejection_channels_314__flag <= 1'b1;
			end else begin
				ejection_channels_314__flag<= 1'b0;
			end
			if(!(ejection_channels_313__gfpga === ejection_channels_313__bench) && !(ejection_channels_313__bench === 1'bx)) begin
				ejection_channels_313__flag <= 1'b1;
			end else begin
				ejection_channels_313__flag<= 1'b0;
			end
			if(!(ejection_channels_312__gfpga === ejection_channels_312__bench) && !(ejection_channels_312__bench === 1'bx)) begin
				ejection_channels_312__flag <= 1'b1;
			end else begin
				ejection_channels_312__flag<= 1'b0;
			end
			if(!(ejection_channels_311__gfpga === ejection_channels_311__bench) && !(ejection_channels_311__bench === 1'bx)) begin
				ejection_channels_311__flag <= 1'b1;
			end else begin
				ejection_channels_311__flag<= 1'b0;
			end
			if(!(ejection_channels_310__gfpga === ejection_channels_310__bench) && !(ejection_channels_310__bench === 1'bx)) begin
				ejection_channels_310__flag <= 1'b1;
			end else begin
				ejection_channels_310__flag<= 1'b0;
			end
			if(!(ejection_channels_309__gfpga === ejection_channels_309__bench) && !(ejection_channels_309__bench === 1'bx)) begin
				ejection_channels_309__flag <= 1'b1;
			end else begin
				ejection_channels_309__flag<= 1'b0;
			end
			if(!(ejection_channels_308__gfpga === ejection_channels_308__bench) && !(ejection_channels_308__bench === 1'bx)) begin
				ejection_channels_308__flag <= 1'b1;
			end else begin
				ejection_channels_308__flag<= 1'b0;
			end
			if(!(ejection_channels_307__gfpga === ejection_channels_307__bench) && !(ejection_channels_307__bench === 1'bx)) begin
				ejection_channels_307__flag <= 1'b1;
			end else begin
				ejection_channels_307__flag<= 1'b0;
			end
			if(!(ejection_channels_306__gfpga === ejection_channels_306__bench) && !(ejection_channels_306__bench === 1'bx)) begin
				ejection_channels_306__flag <= 1'b1;
			end else begin
				ejection_channels_306__flag<= 1'b0;
			end
			if(!(ejection_channels_305__gfpga === ejection_channels_305__bench) && !(ejection_channels_305__bench === 1'bx)) begin
				ejection_channels_305__flag <= 1'b1;
			end else begin
				ejection_channels_305__flag<= 1'b0;
			end
			if(!(ejection_channels_304__gfpga === ejection_channels_304__bench) && !(ejection_channels_304__bench === 1'bx)) begin
				ejection_channels_304__flag <= 1'b1;
			end else begin
				ejection_channels_304__flag<= 1'b0;
			end
			if(!(ejection_channels_303__gfpga === ejection_channels_303__bench) && !(ejection_channels_303__bench === 1'bx)) begin
				ejection_channels_303__flag <= 1'b1;
			end else begin
				ejection_channels_303__flag<= 1'b0;
			end
			if(!(ejection_channels_302__gfpga === ejection_channels_302__bench) && !(ejection_channels_302__bench === 1'bx)) begin
				ejection_channels_302__flag <= 1'b1;
			end else begin
				ejection_channels_302__flag<= 1'b0;
			end
			if(!(ejection_channels_301__gfpga === ejection_channels_301__bench) && !(ejection_channels_301__bench === 1'bx)) begin
				ejection_channels_301__flag <= 1'b1;
			end else begin
				ejection_channels_301__flag<= 1'b0;
			end
			if(!(ejection_channels_300__gfpga === ejection_channels_300__bench) && !(ejection_channels_300__bench === 1'bx)) begin
				ejection_channels_300__flag <= 1'b1;
			end else begin
				ejection_channels_300__flag<= 1'b0;
			end
			if(!(ejection_channels_299__gfpga === ejection_channels_299__bench) && !(ejection_channels_299__bench === 1'bx)) begin
				ejection_channels_299__flag <= 1'b1;
			end else begin
				ejection_channels_299__flag<= 1'b0;
			end
			if(!(ejection_channels_298__gfpga === ejection_channels_298__bench) && !(ejection_channels_298__bench === 1'bx)) begin
				ejection_channels_298__flag <= 1'b1;
			end else begin
				ejection_channels_298__flag<= 1'b0;
			end
			if(!(ejection_channels_297__gfpga === ejection_channels_297__bench) && !(ejection_channels_297__bench === 1'bx)) begin
				ejection_channels_297__flag <= 1'b1;
			end else begin
				ejection_channels_297__flag<= 1'b0;
			end
			if(!(ejection_channels_296__gfpga === ejection_channels_296__bench) && !(ejection_channels_296__bench === 1'bx)) begin
				ejection_channels_296__flag <= 1'b1;
			end else begin
				ejection_channels_296__flag<= 1'b0;
			end
			if(!(ejection_channels_295__gfpga === ejection_channels_295__bench) && !(ejection_channels_295__bench === 1'bx)) begin
				ejection_channels_295__flag <= 1'b1;
			end else begin
				ejection_channels_295__flag<= 1'b0;
			end
			if(!(ejection_channels_294__gfpga === ejection_channels_294__bench) && !(ejection_channels_294__bench === 1'bx)) begin
				ejection_channels_294__flag <= 1'b1;
			end else begin
				ejection_channels_294__flag<= 1'b0;
			end
			if(!(ejection_channels_293__gfpga === ejection_channels_293__bench) && !(ejection_channels_293__bench === 1'bx)) begin
				ejection_channels_293__flag <= 1'b1;
			end else begin
				ejection_channels_293__flag<= 1'b0;
			end
			if(!(ejection_channels_292__gfpga === ejection_channels_292__bench) && !(ejection_channels_292__bench === 1'bx)) begin
				ejection_channels_292__flag <= 1'b1;
			end else begin
				ejection_channels_292__flag<= 1'b0;
			end
			if(!(ejection_channels_291__gfpga === ejection_channels_291__bench) && !(ejection_channels_291__bench === 1'bx)) begin
				ejection_channels_291__flag <= 1'b1;
			end else begin
				ejection_channels_291__flag<= 1'b0;
			end
			if(!(ejection_channels_290__gfpga === ejection_channels_290__bench) && !(ejection_channels_290__bench === 1'bx)) begin
				ejection_channels_290__flag <= 1'b1;
			end else begin
				ejection_channels_290__flag<= 1'b0;
			end
			if(!(ejection_channels_289__gfpga === ejection_channels_289__bench) && !(ejection_channels_289__bench === 1'bx)) begin
				ejection_channels_289__flag <= 1'b1;
			end else begin
				ejection_channels_289__flag<= 1'b0;
			end
			if(!(ejection_channels_288__gfpga === ejection_channels_288__bench) && !(ejection_channels_288__bench === 1'bx)) begin
				ejection_channels_288__flag <= 1'b1;
			end else begin
				ejection_channels_288__flag<= 1'b0;
			end
			if(!(ejection_channels_287__gfpga === ejection_channels_287__bench) && !(ejection_channels_287__bench === 1'bx)) begin
				ejection_channels_287__flag <= 1'b1;
			end else begin
				ejection_channels_287__flag<= 1'b0;
			end
			if(!(ejection_channels_286__gfpga === ejection_channels_286__bench) && !(ejection_channels_286__bench === 1'bx)) begin
				ejection_channels_286__flag <= 1'b1;
			end else begin
				ejection_channels_286__flag<= 1'b0;
			end
			if(!(ejection_channels_285__gfpga === ejection_channels_285__bench) && !(ejection_channels_285__bench === 1'bx)) begin
				ejection_channels_285__flag <= 1'b1;
			end else begin
				ejection_channels_285__flag<= 1'b0;
			end
			if(!(ejection_channels_284__gfpga === ejection_channels_284__bench) && !(ejection_channels_284__bench === 1'bx)) begin
				ejection_channels_284__flag <= 1'b1;
			end else begin
				ejection_channels_284__flag<= 1'b0;
			end
			if(!(ejection_channels_283__gfpga === ejection_channels_283__bench) && !(ejection_channels_283__bench === 1'bx)) begin
				ejection_channels_283__flag <= 1'b1;
			end else begin
				ejection_channels_283__flag<= 1'b0;
			end
			if(!(ejection_channels_282__gfpga === ejection_channels_282__bench) && !(ejection_channels_282__bench === 1'bx)) begin
				ejection_channels_282__flag <= 1'b1;
			end else begin
				ejection_channels_282__flag<= 1'b0;
			end
			if(!(ejection_channels_281__gfpga === ejection_channels_281__bench) && !(ejection_channels_281__bench === 1'bx)) begin
				ejection_channels_281__flag <= 1'b1;
			end else begin
				ejection_channels_281__flag<= 1'b0;
			end
			if(!(ejection_channels_280__gfpga === ejection_channels_280__bench) && !(ejection_channels_280__bench === 1'bx)) begin
				ejection_channels_280__flag <= 1'b1;
			end else begin
				ejection_channels_280__flag<= 1'b0;
			end
			if(!(ejection_channels_279__gfpga === ejection_channels_279__bench) && !(ejection_channels_279__bench === 1'bx)) begin
				ejection_channels_279__flag <= 1'b1;
			end else begin
				ejection_channels_279__flag<= 1'b0;
			end
			if(!(ejection_channels_278__gfpga === ejection_channels_278__bench) && !(ejection_channels_278__bench === 1'bx)) begin
				ejection_channels_278__flag <= 1'b1;
			end else begin
				ejection_channels_278__flag<= 1'b0;
			end
			if(!(ejection_channels_277__gfpga === ejection_channels_277__bench) && !(ejection_channels_277__bench === 1'bx)) begin
				ejection_channels_277__flag <= 1'b1;
			end else begin
				ejection_channels_277__flag<= 1'b0;
			end
			if(!(ejection_channels_276__gfpga === ejection_channels_276__bench) && !(ejection_channels_276__bench === 1'bx)) begin
				ejection_channels_276__flag <= 1'b1;
			end else begin
				ejection_channels_276__flag<= 1'b0;
			end
			if(!(ejection_channels_275__gfpga === ejection_channels_275__bench) && !(ejection_channels_275__bench === 1'bx)) begin
				ejection_channels_275__flag <= 1'b1;
			end else begin
				ejection_channels_275__flag<= 1'b0;
			end
			if(!(ejection_channels_274__gfpga === ejection_channels_274__bench) && !(ejection_channels_274__bench === 1'bx)) begin
				ejection_channels_274__flag <= 1'b1;
			end else begin
				ejection_channels_274__flag<= 1'b0;
			end
			if(!(ejection_channels_273__gfpga === ejection_channels_273__bench) && !(ejection_channels_273__bench === 1'bx)) begin
				ejection_channels_273__flag <= 1'b1;
			end else begin
				ejection_channels_273__flag<= 1'b0;
			end
			if(!(ejection_channels_272__gfpga === ejection_channels_272__bench) && !(ejection_channels_272__bench === 1'bx)) begin
				ejection_channels_272__flag <= 1'b1;
			end else begin
				ejection_channels_272__flag<= 1'b0;
			end
			if(!(ejection_channels_271__gfpga === ejection_channels_271__bench) && !(ejection_channels_271__bench === 1'bx)) begin
				ejection_channels_271__flag <= 1'b1;
			end else begin
				ejection_channels_271__flag<= 1'b0;
			end
			if(!(ejection_channels_270__gfpga === ejection_channels_270__bench) && !(ejection_channels_270__bench === 1'bx)) begin
				ejection_channels_270__flag <= 1'b1;
			end else begin
				ejection_channels_270__flag<= 1'b0;
			end
			if(!(ejection_channels_269__gfpga === ejection_channels_269__bench) && !(ejection_channels_269__bench === 1'bx)) begin
				ejection_channels_269__flag <= 1'b1;
			end else begin
				ejection_channels_269__flag<= 1'b0;
			end
			if(!(ejection_channels_268__gfpga === ejection_channels_268__bench) && !(ejection_channels_268__bench === 1'bx)) begin
				ejection_channels_268__flag <= 1'b1;
			end else begin
				ejection_channels_268__flag<= 1'b0;
			end
			if(!(ejection_channels_267__gfpga === ejection_channels_267__bench) && !(ejection_channels_267__bench === 1'bx)) begin
				ejection_channels_267__flag <= 1'b1;
			end else begin
				ejection_channels_267__flag<= 1'b0;
			end
			if(!(ejection_channels_266__gfpga === ejection_channels_266__bench) && !(ejection_channels_266__bench === 1'bx)) begin
				ejection_channels_266__flag <= 1'b1;
			end else begin
				ejection_channels_266__flag<= 1'b0;
			end
			if(!(ejection_channels_265__gfpga === ejection_channels_265__bench) && !(ejection_channels_265__bench === 1'bx)) begin
				ejection_channels_265__flag <= 1'b1;
			end else begin
				ejection_channels_265__flag<= 1'b0;
			end
			if(!(ejection_channels_264__gfpga === ejection_channels_264__bench) && !(ejection_channels_264__bench === 1'bx)) begin
				ejection_channels_264__flag <= 1'b1;
			end else begin
				ejection_channels_264__flag<= 1'b0;
			end
			if(!(ejection_channels_263__gfpga === ejection_channels_263__bench) && !(ejection_channels_263__bench === 1'bx)) begin
				ejection_channels_263__flag <= 1'b1;
			end else begin
				ejection_channels_263__flag<= 1'b0;
			end
			if(!(ejection_channels_262__gfpga === ejection_channels_262__bench) && !(ejection_channels_262__bench === 1'bx)) begin
				ejection_channels_262__flag <= 1'b1;
			end else begin
				ejection_channels_262__flag<= 1'b0;
			end
			if(!(ejection_channels_261__gfpga === ejection_channels_261__bench) && !(ejection_channels_261__bench === 1'bx)) begin
				ejection_channels_261__flag <= 1'b1;
			end else begin
				ejection_channels_261__flag<= 1'b0;
			end
			if(!(ejection_channels_260__gfpga === ejection_channels_260__bench) && !(ejection_channels_260__bench === 1'bx)) begin
				ejection_channels_260__flag <= 1'b1;
			end else begin
				ejection_channels_260__flag<= 1'b0;
			end
			if(!(ejection_channels_259__gfpga === ejection_channels_259__bench) && !(ejection_channels_259__bench === 1'bx)) begin
				ejection_channels_259__flag <= 1'b1;
			end else begin
				ejection_channels_259__flag<= 1'b0;
			end
			if(!(ejection_channels_258__gfpga === ejection_channels_258__bench) && !(ejection_channels_258__bench === 1'bx)) begin
				ejection_channels_258__flag <= 1'b1;
			end else begin
				ejection_channels_258__flag<= 1'b0;
			end
			if(!(ejection_channels_257__gfpga === ejection_channels_257__bench) && !(ejection_channels_257__bench === 1'bx)) begin
				ejection_channels_257__flag <= 1'b1;
			end else begin
				ejection_channels_257__flag<= 1'b0;
			end
			if(!(ejection_channels_256__gfpga === ejection_channels_256__bench) && !(ejection_channels_256__bench === 1'bx)) begin
				ejection_channels_256__flag <= 1'b1;
			end else begin
				ejection_channels_256__flag<= 1'b0;
			end
			if(!(ejection_channels_255__gfpga === ejection_channels_255__bench) && !(ejection_channels_255__bench === 1'bx)) begin
				ejection_channels_255__flag <= 1'b1;
			end else begin
				ejection_channels_255__flag<= 1'b0;
			end
			if(!(ejection_channels_254__gfpga === ejection_channels_254__bench) && !(ejection_channels_254__bench === 1'bx)) begin
				ejection_channels_254__flag <= 1'b1;
			end else begin
				ejection_channels_254__flag<= 1'b0;
			end
			if(!(ejection_channels_253__gfpga === ejection_channels_253__bench) && !(ejection_channels_253__bench === 1'bx)) begin
				ejection_channels_253__flag <= 1'b1;
			end else begin
				ejection_channels_253__flag<= 1'b0;
			end
			if(!(ejection_channels_252__gfpga === ejection_channels_252__bench) && !(ejection_channels_252__bench === 1'bx)) begin
				ejection_channels_252__flag <= 1'b1;
			end else begin
				ejection_channels_252__flag<= 1'b0;
			end
			if(!(ejection_channels_251__gfpga === ejection_channels_251__bench) && !(ejection_channels_251__bench === 1'bx)) begin
				ejection_channels_251__flag <= 1'b1;
			end else begin
				ejection_channels_251__flag<= 1'b0;
			end
			if(!(ejection_channels_250__gfpga === ejection_channels_250__bench) && !(ejection_channels_250__bench === 1'bx)) begin
				ejection_channels_250__flag <= 1'b1;
			end else begin
				ejection_channels_250__flag<= 1'b0;
			end
			if(!(ejection_channels_249__gfpga === ejection_channels_249__bench) && !(ejection_channels_249__bench === 1'bx)) begin
				ejection_channels_249__flag <= 1'b1;
			end else begin
				ejection_channels_249__flag<= 1'b0;
			end
			if(!(ejection_channels_248__gfpga === ejection_channels_248__bench) && !(ejection_channels_248__bench === 1'bx)) begin
				ejection_channels_248__flag <= 1'b1;
			end else begin
				ejection_channels_248__flag<= 1'b0;
			end
			if(!(ejection_channels_247__gfpga === ejection_channels_247__bench) && !(ejection_channels_247__bench === 1'bx)) begin
				ejection_channels_247__flag <= 1'b1;
			end else begin
				ejection_channels_247__flag<= 1'b0;
			end
			if(!(ejection_channels_246__gfpga === ejection_channels_246__bench) && !(ejection_channels_246__bench === 1'bx)) begin
				ejection_channels_246__flag <= 1'b1;
			end else begin
				ejection_channels_246__flag<= 1'b0;
			end
			if(!(ejection_channels_245__gfpga === ejection_channels_245__bench) && !(ejection_channels_245__bench === 1'bx)) begin
				ejection_channels_245__flag <= 1'b1;
			end else begin
				ejection_channels_245__flag<= 1'b0;
			end
			if(!(ejection_channels_244__gfpga === ejection_channels_244__bench) && !(ejection_channels_244__bench === 1'bx)) begin
				ejection_channels_244__flag <= 1'b1;
			end else begin
				ejection_channels_244__flag<= 1'b0;
			end
			if(!(ejection_channels_243__gfpga === ejection_channels_243__bench) && !(ejection_channels_243__bench === 1'bx)) begin
				ejection_channels_243__flag <= 1'b1;
			end else begin
				ejection_channels_243__flag<= 1'b0;
			end
			if(!(ejection_channels_242__gfpga === ejection_channels_242__bench) && !(ejection_channels_242__bench === 1'bx)) begin
				ejection_channels_242__flag <= 1'b1;
			end else begin
				ejection_channels_242__flag<= 1'b0;
			end
			if(!(ejection_channels_241__gfpga === ejection_channels_241__bench) && !(ejection_channels_241__bench === 1'bx)) begin
				ejection_channels_241__flag <= 1'b1;
			end else begin
				ejection_channels_241__flag<= 1'b0;
			end
			if(!(ejection_channels_240__gfpga === ejection_channels_240__bench) && !(ejection_channels_240__bench === 1'bx)) begin
				ejection_channels_240__flag <= 1'b1;
			end else begin
				ejection_channels_240__flag<= 1'b0;
			end
			if(!(ejection_channels_239__gfpga === ejection_channels_239__bench) && !(ejection_channels_239__bench === 1'bx)) begin
				ejection_channels_239__flag <= 1'b1;
			end else begin
				ejection_channels_239__flag<= 1'b0;
			end
			if(!(ejection_channels_238__gfpga === ejection_channels_238__bench) && !(ejection_channels_238__bench === 1'bx)) begin
				ejection_channels_238__flag <= 1'b1;
			end else begin
				ejection_channels_238__flag<= 1'b0;
			end
			if(!(ejection_channels_237__gfpga === ejection_channels_237__bench) && !(ejection_channels_237__bench === 1'bx)) begin
				ejection_channels_237__flag <= 1'b1;
			end else begin
				ejection_channels_237__flag<= 1'b0;
			end
			if(!(ejection_channels_236__gfpga === ejection_channels_236__bench) && !(ejection_channels_236__bench === 1'bx)) begin
				ejection_channels_236__flag <= 1'b1;
			end else begin
				ejection_channels_236__flag<= 1'b0;
			end
			if(!(ejection_channels_235__gfpga === ejection_channels_235__bench) && !(ejection_channels_235__bench === 1'bx)) begin
				ejection_channels_235__flag <= 1'b1;
			end else begin
				ejection_channels_235__flag<= 1'b0;
			end
			if(!(ejection_channels_234__gfpga === ejection_channels_234__bench) && !(ejection_channels_234__bench === 1'bx)) begin
				ejection_channels_234__flag <= 1'b1;
			end else begin
				ejection_channels_234__flag<= 1'b0;
			end
			if(!(ejection_channels_233__gfpga === ejection_channels_233__bench) && !(ejection_channels_233__bench === 1'bx)) begin
				ejection_channels_233__flag <= 1'b1;
			end else begin
				ejection_channels_233__flag<= 1'b0;
			end
			if(!(ejection_channels_232__gfpga === ejection_channels_232__bench) && !(ejection_channels_232__bench === 1'bx)) begin
				ejection_channels_232__flag <= 1'b1;
			end else begin
				ejection_channels_232__flag<= 1'b0;
			end
			if(!(ejection_channels_231__gfpga === ejection_channels_231__bench) && !(ejection_channels_231__bench === 1'bx)) begin
				ejection_channels_231__flag <= 1'b1;
			end else begin
				ejection_channels_231__flag<= 1'b0;
			end
			if(!(ejection_channels_230__gfpga === ejection_channels_230__bench) && !(ejection_channels_230__bench === 1'bx)) begin
				ejection_channels_230__flag <= 1'b1;
			end else begin
				ejection_channels_230__flag<= 1'b0;
			end
			if(!(ejection_channels_229__gfpga === ejection_channels_229__bench) && !(ejection_channels_229__bench === 1'bx)) begin
				ejection_channels_229__flag <= 1'b1;
			end else begin
				ejection_channels_229__flag<= 1'b0;
			end
			if(!(ejection_channels_228__gfpga === ejection_channels_228__bench) && !(ejection_channels_228__bench === 1'bx)) begin
				ejection_channels_228__flag <= 1'b1;
			end else begin
				ejection_channels_228__flag<= 1'b0;
			end
			if(!(ejection_channels_227__gfpga === ejection_channels_227__bench) && !(ejection_channels_227__bench === 1'bx)) begin
				ejection_channels_227__flag <= 1'b1;
			end else begin
				ejection_channels_227__flag<= 1'b0;
			end
			if(!(ejection_channels_226__gfpga === ejection_channels_226__bench) && !(ejection_channels_226__bench === 1'bx)) begin
				ejection_channels_226__flag <= 1'b1;
			end else begin
				ejection_channels_226__flag<= 1'b0;
			end
			if(!(ejection_channels_225__gfpga === ejection_channels_225__bench) && !(ejection_channels_225__bench === 1'bx)) begin
				ejection_channels_225__flag <= 1'b1;
			end else begin
				ejection_channels_225__flag<= 1'b0;
			end
			if(!(ejection_channels_224__gfpga === ejection_channels_224__bench) && !(ejection_channels_224__bench === 1'bx)) begin
				ejection_channels_224__flag <= 1'b1;
			end else begin
				ejection_channels_224__flag<= 1'b0;
			end
			if(!(ejection_channels_223__gfpga === ejection_channels_223__bench) && !(ejection_channels_223__bench === 1'bx)) begin
				ejection_channels_223__flag <= 1'b1;
			end else begin
				ejection_channels_223__flag<= 1'b0;
			end
			if(!(ejection_channels_222__gfpga === ejection_channels_222__bench) && !(ejection_channels_222__bench === 1'bx)) begin
				ejection_channels_222__flag <= 1'b1;
			end else begin
				ejection_channels_222__flag<= 1'b0;
			end
			if(!(ejection_channels_221__gfpga === ejection_channels_221__bench) && !(ejection_channels_221__bench === 1'bx)) begin
				ejection_channels_221__flag <= 1'b1;
			end else begin
				ejection_channels_221__flag<= 1'b0;
			end
			if(!(ejection_channels_220__gfpga === ejection_channels_220__bench) && !(ejection_channels_220__bench === 1'bx)) begin
				ejection_channels_220__flag <= 1'b1;
			end else begin
				ejection_channels_220__flag<= 1'b0;
			end
			if(!(ejection_channels_219__gfpga === ejection_channels_219__bench) && !(ejection_channels_219__bench === 1'bx)) begin
				ejection_channels_219__flag <= 1'b1;
			end else begin
				ejection_channels_219__flag<= 1'b0;
			end
			if(!(ejection_channels_218__gfpga === ejection_channels_218__bench) && !(ejection_channels_218__bench === 1'bx)) begin
				ejection_channels_218__flag <= 1'b1;
			end else begin
				ejection_channels_218__flag<= 1'b0;
			end
			if(!(ejection_channels_217__gfpga === ejection_channels_217__bench) && !(ejection_channels_217__bench === 1'bx)) begin
				ejection_channels_217__flag <= 1'b1;
			end else begin
				ejection_channels_217__flag<= 1'b0;
			end
			if(!(ejection_channels_216__gfpga === ejection_channels_216__bench) && !(ejection_channels_216__bench === 1'bx)) begin
				ejection_channels_216__flag <= 1'b1;
			end else begin
				ejection_channels_216__flag<= 1'b0;
			end
			if(!(ejection_channels_215__gfpga === ejection_channels_215__bench) && !(ejection_channels_215__bench === 1'bx)) begin
				ejection_channels_215__flag <= 1'b1;
			end else begin
				ejection_channels_215__flag<= 1'b0;
			end
			if(!(ejection_channels_214__gfpga === ejection_channels_214__bench) && !(ejection_channels_214__bench === 1'bx)) begin
				ejection_channels_214__flag <= 1'b1;
			end else begin
				ejection_channels_214__flag<= 1'b0;
			end
			if(!(ejection_channels_213__gfpga === ejection_channels_213__bench) && !(ejection_channels_213__bench === 1'bx)) begin
				ejection_channels_213__flag <= 1'b1;
			end else begin
				ejection_channels_213__flag<= 1'b0;
			end
			if(!(ejection_channels_212__gfpga === ejection_channels_212__bench) && !(ejection_channels_212__bench === 1'bx)) begin
				ejection_channels_212__flag <= 1'b1;
			end else begin
				ejection_channels_212__flag<= 1'b0;
			end
			if(!(ejection_channels_211__gfpga === ejection_channels_211__bench) && !(ejection_channels_211__bench === 1'bx)) begin
				ejection_channels_211__flag <= 1'b1;
			end else begin
				ejection_channels_211__flag<= 1'b0;
			end
			if(!(ejection_channels_210__gfpga === ejection_channels_210__bench) && !(ejection_channels_210__bench === 1'bx)) begin
				ejection_channels_210__flag <= 1'b1;
			end else begin
				ejection_channels_210__flag<= 1'b0;
			end
			if(!(ejection_channels_209__gfpga === ejection_channels_209__bench) && !(ejection_channels_209__bench === 1'bx)) begin
				ejection_channels_209__flag <= 1'b1;
			end else begin
				ejection_channels_209__flag<= 1'b0;
			end
			if(!(ejection_channels_208__gfpga === ejection_channels_208__bench) && !(ejection_channels_208__bench === 1'bx)) begin
				ejection_channels_208__flag <= 1'b1;
			end else begin
				ejection_channels_208__flag<= 1'b0;
			end
			if(!(ejection_channels_207__gfpga === ejection_channels_207__bench) && !(ejection_channels_207__bench === 1'bx)) begin
				ejection_channels_207__flag <= 1'b1;
			end else begin
				ejection_channels_207__flag<= 1'b0;
			end
			if(!(ejection_channels_206__gfpga === ejection_channels_206__bench) && !(ejection_channels_206__bench === 1'bx)) begin
				ejection_channels_206__flag <= 1'b1;
			end else begin
				ejection_channels_206__flag<= 1'b0;
			end
			if(!(ejection_channels_205__gfpga === ejection_channels_205__bench) && !(ejection_channels_205__bench === 1'bx)) begin
				ejection_channels_205__flag <= 1'b1;
			end else begin
				ejection_channels_205__flag<= 1'b0;
			end
			if(!(ejection_channels_204__gfpga === ejection_channels_204__bench) && !(ejection_channels_204__bench === 1'bx)) begin
				ejection_channels_204__flag <= 1'b1;
			end else begin
				ejection_channels_204__flag<= 1'b0;
			end
			if(!(ejection_channels_203__gfpga === ejection_channels_203__bench) && !(ejection_channels_203__bench === 1'bx)) begin
				ejection_channels_203__flag <= 1'b1;
			end else begin
				ejection_channels_203__flag<= 1'b0;
			end
			if(!(ejection_channels_202__gfpga === ejection_channels_202__bench) && !(ejection_channels_202__bench === 1'bx)) begin
				ejection_channels_202__flag <= 1'b1;
			end else begin
				ejection_channels_202__flag<= 1'b0;
			end
			if(!(ejection_channels_201__gfpga === ejection_channels_201__bench) && !(ejection_channels_201__bench === 1'bx)) begin
				ejection_channels_201__flag <= 1'b1;
			end else begin
				ejection_channels_201__flag<= 1'b0;
			end
			if(!(ejection_channels_200__gfpga === ejection_channels_200__bench) && !(ejection_channels_200__bench === 1'bx)) begin
				ejection_channels_200__flag <= 1'b1;
			end else begin
				ejection_channels_200__flag<= 1'b0;
			end
			if(!(ejection_channels_199__gfpga === ejection_channels_199__bench) && !(ejection_channels_199__bench === 1'bx)) begin
				ejection_channels_199__flag <= 1'b1;
			end else begin
				ejection_channels_199__flag<= 1'b0;
			end
			if(!(ejection_channels_198__gfpga === ejection_channels_198__bench) && !(ejection_channels_198__bench === 1'bx)) begin
				ejection_channels_198__flag <= 1'b1;
			end else begin
				ejection_channels_198__flag<= 1'b0;
			end
			if(!(ejection_channels_197__gfpga === ejection_channels_197__bench) && !(ejection_channels_197__bench === 1'bx)) begin
				ejection_channels_197__flag <= 1'b1;
			end else begin
				ejection_channels_197__flag<= 1'b0;
			end
			if(!(ejection_channels_196__gfpga === ejection_channels_196__bench) && !(ejection_channels_196__bench === 1'bx)) begin
				ejection_channels_196__flag <= 1'b1;
			end else begin
				ejection_channels_196__flag<= 1'b0;
			end
			if(!(ejection_channels_195__gfpga === ejection_channels_195__bench) && !(ejection_channels_195__bench === 1'bx)) begin
				ejection_channels_195__flag <= 1'b1;
			end else begin
				ejection_channels_195__flag<= 1'b0;
			end
			if(!(ejection_channels_194__gfpga === ejection_channels_194__bench) && !(ejection_channels_194__bench === 1'bx)) begin
				ejection_channels_194__flag <= 1'b1;
			end else begin
				ejection_channels_194__flag<= 1'b0;
			end
			if(!(ejection_channels_193__gfpga === ejection_channels_193__bench) && !(ejection_channels_193__bench === 1'bx)) begin
				ejection_channels_193__flag <= 1'b1;
			end else begin
				ejection_channels_193__flag<= 1'b0;
			end
			if(!(ejection_channels_192__gfpga === ejection_channels_192__bench) && !(ejection_channels_192__bench === 1'bx)) begin
				ejection_channels_192__flag <= 1'b1;
			end else begin
				ejection_channels_192__flag<= 1'b0;
			end
			if(!(ejection_channels_191__gfpga === ejection_channels_191__bench) && !(ejection_channels_191__bench === 1'bx)) begin
				ejection_channels_191__flag <= 1'b1;
			end else begin
				ejection_channels_191__flag<= 1'b0;
			end
			if(!(ejection_channels_190__gfpga === ejection_channels_190__bench) && !(ejection_channels_190__bench === 1'bx)) begin
				ejection_channels_190__flag <= 1'b1;
			end else begin
				ejection_channels_190__flag<= 1'b0;
			end
			if(!(ejection_channels_189__gfpga === ejection_channels_189__bench) && !(ejection_channels_189__bench === 1'bx)) begin
				ejection_channels_189__flag <= 1'b1;
			end else begin
				ejection_channels_189__flag<= 1'b0;
			end
			if(!(ejection_channels_188__gfpga === ejection_channels_188__bench) && !(ejection_channels_188__bench === 1'bx)) begin
				ejection_channels_188__flag <= 1'b1;
			end else begin
				ejection_channels_188__flag<= 1'b0;
			end
			if(!(ejection_channels_187__gfpga === ejection_channels_187__bench) && !(ejection_channels_187__bench === 1'bx)) begin
				ejection_channels_187__flag <= 1'b1;
			end else begin
				ejection_channels_187__flag<= 1'b0;
			end
			if(!(ejection_channels_186__gfpga === ejection_channels_186__bench) && !(ejection_channels_186__bench === 1'bx)) begin
				ejection_channels_186__flag <= 1'b1;
			end else begin
				ejection_channels_186__flag<= 1'b0;
			end
			if(!(ejection_channels_185__gfpga === ejection_channels_185__bench) && !(ejection_channels_185__bench === 1'bx)) begin
				ejection_channels_185__flag <= 1'b1;
			end else begin
				ejection_channels_185__flag<= 1'b0;
			end
			if(!(ejection_channels_184__gfpga === ejection_channels_184__bench) && !(ejection_channels_184__bench === 1'bx)) begin
				ejection_channels_184__flag <= 1'b1;
			end else begin
				ejection_channels_184__flag<= 1'b0;
			end
			if(!(ejection_channels_183__gfpga === ejection_channels_183__bench) && !(ejection_channels_183__bench === 1'bx)) begin
				ejection_channels_183__flag <= 1'b1;
			end else begin
				ejection_channels_183__flag<= 1'b0;
			end
			if(!(ejection_channels_182__gfpga === ejection_channels_182__bench) && !(ejection_channels_182__bench === 1'bx)) begin
				ejection_channels_182__flag <= 1'b1;
			end else begin
				ejection_channels_182__flag<= 1'b0;
			end
			if(!(ejection_channels_181__gfpga === ejection_channels_181__bench) && !(ejection_channels_181__bench === 1'bx)) begin
				ejection_channels_181__flag <= 1'b1;
			end else begin
				ejection_channels_181__flag<= 1'b0;
			end
			if(!(ejection_channels_180__gfpga === ejection_channels_180__bench) && !(ejection_channels_180__bench === 1'bx)) begin
				ejection_channels_180__flag <= 1'b1;
			end else begin
				ejection_channels_180__flag<= 1'b0;
			end
			if(!(ejection_channels_179__gfpga === ejection_channels_179__bench) && !(ejection_channels_179__bench === 1'bx)) begin
				ejection_channels_179__flag <= 1'b1;
			end else begin
				ejection_channels_179__flag<= 1'b0;
			end
			if(!(ejection_channels_178__gfpga === ejection_channels_178__bench) && !(ejection_channels_178__bench === 1'bx)) begin
				ejection_channels_178__flag <= 1'b1;
			end else begin
				ejection_channels_178__flag<= 1'b0;
			end
			if(!(ejection_channels_177__gfpga === ejection_channels_177__bench) && !(ejection_channels_177__bench === 1'bx)) begin
				ejection_channels_177__flag <= 1'b1;
			end else begin
				ejection_channels_177__flag<= 1'b0;
			end
			if(!(ejection_channels_176__gfpga === ejection_channels_176__bench) && !(ejection_channels_176__bench === 1'bx)) begin
				ejection_channels_176__flag <= 1'b1;
			end else begin
				ejection_channels_176__flag<= 1'b0;
			end
			if(!(ejection_channels_175__gfpga === ejection_channels_175__bench) && !(ejection_channels_175__bench === 1'bx)) begin
				ejection_channels_175__flag <= 1'b1;
			end else begin
				ejection_channels_175__flag<= 1'b0;
			end
			if(!(ejection_channels_174__gfpga === ejection_channels_174__bench) && !(ejection_channels_174__bench === 1'bx)) begin
				ejection_channels_174__flag <= 1'b1;
			end else begin
				ejection_channels_174__flag<= 1'b0;
			end
			if(!(ejection_channels_173__gfpga === ejection_channels_173__bench) && !(ejection_channels_173__bench === 1'bx)) begin
				ejection_channels_173__flag <= 1'b1;
			end else begin
				ejection_channels_173__flag<= 1'b0;
			end
			if(!(ejection_channels_172__gfpga === ejection_channels_172__bench) && !(ejection_channels_172__bench === 1'bx)) begin
				ejection_channels_172__flag <= 1'b1;
			end else begin
				ejection_channels_172__flag<= 1'b0;
			end
			if(!(ejection_channels_171__gfpga === ejection_channels_171__bench) && !(ejection_channels_171__bench === 1'bx)) begin
				ejection_channels_171__flag <= 1'b1;
			end else begin
				ejection_channels_171__flag<= 1'b0;
			end
			if(!(ejection_channels_170__gfpga === ejection_channels_170__bench) && !(ejection_channels_170__bench === 1'bx)) begin
				ejection_channels_170__flag <= 1'b1;
			end else begin
				ejection_channels_170__flag<= 1'b0;
			end
			if(!(ejection_channels_169__gfpga === ejection_channels_169__bench) && !(ejection_channels_169__bench === 1'bx)) begin
				ejection_channels_169__flag <= 1'b1;
			end else begin
				ejection_channels_169__flag<= 1'b0;
			end
			if(!(ejection_channels_168__gfpga === ejection_channels_168__bench) && !(ejection_channels_168__bench === 1'bx)) begin
				ejection_channels_168__flag <= 1'b1;
			end else begin
				ejection_channels_168__flag<= 1'b0;
			end
			if(!(ejection_channels_167__gfpga === ejection_channels_167__bench) && !(ejection_channels_167__bench === 1'bx)) begin
				ejection_channels_167__flag <= 1'b1;
			end else begin
				ejection_channels_167__flag<= 1'b0;
			end
			if(!(ejection_channels_166__gfpga === ejection_channels_166__bench) && !(ejection_channels_166__bench === 1'bx)) begin
				ejection_channels_166__flag <= 1'b1;
			end else begin
				ejection_channels_166__flag<= 1'b0;
			end
			if(!(ejection_channels_165__gfpga === ejection_channels_165__bench) && !(ejection_channels_165__bench === 1'bx)) begin
				ejection_channels_165__flag <= 1'b1;
			end else begin
				ejection_channels_165__flag<= 1'b0;
			end
			if(!(ejection_channels_164__gfpga === ejection_channels_164__bench) && !(ejection_channels_164__bench === 1'bx)) begin
				ejection_channels_164__flag <= 1'b1;
			end else begin
				ejection_channels_164__flag<= 1'b0;
			end
			if(!(ejection_channels_163__gfpga === ejection_channels_163__bench) && !(ejection_channels_163__bench === 1'bx)) begin
				ejection_channels_163__flag <= 1'b1;
			end else begin
				ejection_channels_163__flag<= 1'b0;
			end
			if(!(ejection_channels_162__gfpga === ejection_channels_162__bench) && !(ejection_channels_162__bench === 1'bx)) begin
				ejection_channels_162__flag <= 1'b1;
			end else begin
				ejection_channels_162__flag<= 1'b0;
			end
			if(!(ejection_channels_161__gfpga === ejection_channels_161__bench) && !(ejection_channels_161__bench === 1'bx)) begin
				ejection_channels_161__flag <= 1'b1;
			end else begin
				ejection_channels_161__flag<= 1'b0;
			end
			if(!(ejection_channels_160__gfpga === ejection_channels_160__bench) && !(ejection_channels_160__bench === 1'bx)) begin
				ejection_channels_160__flag <= 1'b1;
			end else begin
				ejection_channels_160__flag<= 1'b0;
			end
			if(!(ejection_channels_159__gfpga === ejection_channels_159__bench) && !(ejection_channels_159__bench === 1'bx)) begin
				ejection_channels_159__flag <= 1'b1;
			end else begin
				ejection_channels_159__flag<= 1'b0;
			end
			if(!(ejection_channels_158__gfpga === ejection_channels_158__bench) && !(ejection_channels_158__bench === 1'bx)) begin
				ejection_channels_158__flag <= 1'b1;
			end else begin
				ejection_channels_158__flag<= 1'b0;
			end
			if(!(ejection_channels_157__gfpga === ejection_channels_157__bench) && !(ejection_channels_157__bench === 1'bx)) begin
				ejection_channels_157__flag <= 1'b1;
			end else begin
				ejection_channels_157__flag<= 1'b0;
			end
			if(!(ejection_channels_156__gfpga === ejection_channels_156__bench) && !(ejection_channels_156__bench === 1'bx)) begin
				ejection_channels_156__flag <= 1'b1;
			end else begin
				ejection_channels_156__flag<= 1'b0;
			end
			if(!(ejection_channels_155__gfpga === ejection_channels_155__bench) && !(ejection_channels_155__bench === 1'bx)) begin
				ejection_channels_155__flag <= 1'b1;
			end else begin
				ejection_channels_155__flag<= 1'b0;
			end
			if(!(ejection_channels_154__gfpga === ejection_channels_154__bench) && !(ejection_channels_154__bench === 1'bx)) begin
				ejection_channels_154__flag <= 1'b1;
			end else begin
				ejection_channels_154__flag<= 1'b0;
			end
			if(!(ejection_channels_153__gfpga === ejection_channels_153__bench) && !(ejection_channels_153__bench === 1'bx)) begin
				ejection_channels_153__flag <= 1'b1;
			end else begin
				ejection_channels_153__flag<= 1'b0;
			end
			if(!(ejection_channels_152__gfpga === ejection_channels_152__bench) && !(ejection_channels_152__bench === 1'bx)) begin
				ejection_channels_152__flag <= 1'b1;
			end else begin
				ejection_channels_152__flag<= 1'b0;
			end
			if(!(ejection_channels_151__gfpga === ejection_channels_151__bench) && !(ejection_channels_151__bench === 1'bx)) begin
				ejection_channels_151__flag <= 1'b1;
			end else begin
				ejection_channels_151__flag<= 1'b0;
			end
			if(!(ejection_channels_150__gfpga === ejection_channels_150__bench) && !(ejection_channels_150__bench === 1'bx)) begin
				ejection_channels_150__flag <= 1'b1;
			end else begin
				ejection_channels_150__flag<= 1'b0;
			end
			if(!(ejection_channels_149__gfpga === ejection_channels_149__bench) && !(ejection_channels_149__bench === 1'bx)) begin
				ejection_channels_149__flag <= 1'b1;
			end else begin
				ejection_channels_149__flag<= 1'b0;
			end
			if(!(ejection_channels_148__gfpga === ejection_channels_148__bench) && !(ejection_channels_148__bench === 1'bx)) begin
				ejection_channels_148__flag <= 1'b1;
			end else begin
				ejection_channels_148__flag<= 1'b0;
			end
			if(!(ejection_channels_147__gfpga === ejection_channels_147__bench) && !(ejection_channels_147__bench === 1'bx)) begin
				ejection_channels_147__flag <= 1'b1;
			end else begin
				ejection_channels_147__flag<= 1'b0;
			end
			if(!(ejection_channels_146__gfpga === ejection_channels_146__bench) && !(ejection_channels_146__bench === 1'bx)) begin
				ejection_channels_146__flag <= 1'b1;
			end else begin
				ejection_channels_146__flag<= 1'b0;
			end
			if(!(ejection_channels_145__gfpga === ejection_channels_145__bench) && !(ejection_channels_145__bench === 1'bx)) begin
				ejection_channels_145__flag <= 1'b1;
			end else begin
				ejection_channels_145__flag<= 1'b0;
			end
			if(!(ejection_channels_144__gfpga === ejection_channels_144__bench) && !(ejection_channels_144__bench === 1'bx)) begin
				ejection_channels_144__flag <= 1'b1;
			end else begin
				ejection_channels_144__flag<= 1'b0;
			end
			if(!(ejection_channels_143__gfpga === ejection_channels_143__bench) && !(ejection_channels_143__bench === 1'bx)) begin
				ejection_channels_143__flag <= 1'b1;
			end else begin
				ejection_channels_143__flag<= 1'b0;
			end
			if(!(ejection_channels_142__gfpga === ejection_channels_142__bench) && !(ejection_channels_142__bench === 1'bx)) begin
				ejection_channels_142__flag <= 1'b1;
			end else begin
				ejection_channels_142__flag<= 1'b0;
			end
			if(!(ejection_channels_141__gfpga === ejection_channels_141__bench) && !(ejection_channels_141__bench === 1'bx)) begin
				ejection_channels_141__flag <= 1'b1;
			end else begin
				ejection_channels_141__flag<= 1'b0;
			end
			if(!(ejection_channels_140__gfpga === ejection_channels_140__bench) && !(ejection_channels_140__bench === 1'bx)) begin
				ejection_channels_140__flag <= 1'b1;
			end else begin
				ejection_channels_140__flag<= 1'b0;
			end
			if(!(ejection_channels_139__gfpga === ejection_channels_139__bench) && !(ejection_channels_139__bench === 1'bx)) begin
				ejection_channels_139__flag <= 1'b1;
			end else begin
				ejection_channels_139__flag<= 1'b0;
			end
			if(!(ejection_channels_138__gfpga === ejection_channels_138__bench) && !(ejection_channels_138__bench === 1'bx)) begin
				ejection_channels_138__flag <= 1'b1;
			end else begin
				ejection_channels_138__flag<= 1'b0;
			end
			if(!(ejection_channels_137__gfpga === ejection_channels_137__bench) && !(ejection_channels_137__bench === 1'bx)) begin
				ejection_channels_137__flag <= 1'b1;
			end else begin
				ejection_channels_137__flag<= 1'b0;
			end
			if(!(ejection_channels_136__gfpga === ejection_channels_136__bench) && !(ejection_channels_136__bench === 1'bx)) begin
				ejection_channels_136__flag <= 1'b1;
			end else begin
				ejection_channels_136__flag<= 1'b0;
			end
			if(!(ejection_channels_135__gfpga === ejection_channels_135__bench) && !(ejection_channels_135__bench === 1'bx)) begin
				ejection_channels_135__flag <= 1'b1;
			end else begin
				ejection_channels_135__flag<= 1'b0;
			end
			if(!(ejection_channels_134__gfpga === ejection_channels_134__bench) && !(ejection_channels_134__bench === 1'bx)) begin
				ejection_channels_134__flag <= 1'b1;
			end else begin
				ejection_channels_134__flag<= 1'b0;
			end
			if(!(ejection_channels_133__gfpga === ejection_channels_133__bench) && !(ejection_channels_133__bench === 1'bx)) begin
				ejection_channels_133__flag <= 1'b1;
			end else begin
				ejection_channels_133__flag<= 1'b0;
			end
			if(!(ejection_channels_132__gfpga === ejection_channels_132__bench) && !(ejection_channels_132__bench === 1'bx)) begin
				ejection_channels_132__flag <= 1'b1;
			end else begin
				ejection_channels_132__flag<= 1'b0;
			end
			if(!(ejection_channels_131__gfpga === ejection_channels_131__bench) && !(ejection_channels_131__bench === 1'bx)) begin
				ejection_channels_131__flag <= 1'b1;
			end else begin
				ejection_channels_131__flag<= 1'b0;
			end
			if(!(ejection_channels_130__gfpga === ejection_channels_130__bench) && !(ejection_channels_130__bench === 1'bx)) begin
				ejection_channels_130__flag <= 1'b1;
			end else begin
				ejection_channels_130__flag<= 1'b0;
			end
			if(!(ejection_channels_129__gfpga === ejection_channels_129__bench) && !(ejection_channels_129__bench === 1'bx)) begin
				ejection_channels_129__flag <= 1'b1;
			end else begin
				ejection_channels_129__flag<= 1'b0;
			end
			if(!(ejection_channels_128__gfpga === ejection_channels_128__bench) && !(ejection_channels_128__bench === 1'bx)) begin
				ejection_channels_128__flag <= 1'b1;
			end else begin
				ejection_channels_128__flag<= 1'b0;
			end
			if(!(ejection_channels_127__gfpga === ejection_channels_127__bench) && !(ejection_channels_127__bench === 1'bx)) begin
				ejection_channels_127__flag <= 1'b1;
			end else begin
				ejection_channels_127__flag<= 1'b0;
			end
			if(!(ejection_channels_126__gfpga === ejection_channels_126__bench) && !(ejection_channels_126__bench === 1'bx)) begin
				ejection_channels_126__flag <= 1'b1;
			end else begin
				ejection_channels_126__flag<= 1'b0;
			end
			if(!(ejection_channels_125__gfpga === ejection_channels_125__bench) && !(ejection_channels_125__bench === 1'bx)) begin
				ejection_channels_125__flag <= 1'b1;
			end else begin
				ejection_channels_125__flag<= 1'b0;
			end
			if(!(ejection_channels_124__gfpga === ejection_channels_124__bench) && !(ejection_channels_124__bench === 1'bx)) begin
				ejection_channels_124__flag <= 1'b1;
			end else begin
				ejection_channels_124__flag<= 1'b0;
			end
			if(!(ejection_channels_123__gfpga === ejection_channels_123__bench) && !(ejection_channels_123__bench === 1'bx)) begin
				ejection_channels_123__flag <= 1'b1;
			end else begin
				ejection_channels_123__flag<= 1'b0;
			end
			if(!(ejection_channels_122__gfpga === ejection_channels_122__bench) && !(ejection_channels_122__bench === 1'bx)) begin
				ejection_channels_122__flag <= 1'b1;
			end else begin
				ejection_channels_122__flag<= 1'b0;
			end
			if(!(ejection_channels_121__gfpga === ejection_channels_121__bench) && !(ejection_channels_121__bench === 1'bx)) begin
				ejection_channels_121__flag <= 1'b1;
			end else begin
				ejection_channels_121__flag<= 1'b0;
			end
			if(!(ejection_channels_120__gfpga === ejection_channels_120__bench) && !(ejection_channels_120__bench === 1'bx)) begin
				ejection_channels_120__flag <= 1'b1;
			end else begin
				ejection_channels_120__flag<= 1'b0;
			end
			if(!(ejection_channels_119__gfpga === ejection_channels_119__bench) && !(ejection_channels_119__bench === 1'bx)) begin
				ejection_channels_119__flag <= 1'b1;
			end else begin
				ejection_channels_119__flag<= 1'b0;
			end
			if(!(ejection_channels_118__gfpga === ejection_channels_118__bench) && !(ejection_channels_118__bench === 1'bx)) begin
				ejection_channels_118__flag <= 1'b1;
			end else begin
				ejection_channels_118__flag<= 1'b0;
			end
			if(!(ejection_channels_117__gfpga === ejection_channels_117__bench) && !(ejection_channels_117__bench === 1'bx)) begin
				ejection_channels_117__flag <= 1'b1;
			end else begin
				ejection_channels_117__flag<= 1'b0;
			end
			if(!(ejection_channels_116__gfpga === ejection_channels_116__bench) && !(ejection_channels_116__bench === 1'bx)) begin
				ejection_channels_116__flag <= 1'b1;
			end else begin
				ejection_channels_116__flag<= 1'b0;
			end
			if(!(ejection_channels_115__gfpga === ejection_channels_115__bench) && !(ejection_channels_115__bench === 1'bx)) begin
				ejection_channels_115__flag <= 1'b1;
			end else begin
				ejection_channels_115__flag<= 1'b0;
			end
			if(!(ejection_channels_114__gfpga === ejection_channels_114__bench) && !(ejection_channels_114__bench === 1'bx)) begin
				ejection_channels_114__flag <= 1'b1;
			end else begin
				ejection_channels_114__flag<= 1'b0;
			end
			if(!(ejection_channels_113__gfpga === ejection_channels_113__bench) && !(ejection_channels_113__bench === 1'bx)) begin
				ejection_channels_113__flag <= 1'b1;
			end else begin
				ejection_channels_113__flag<= 1'b0;
			end
			if(!(ejection_channels_112__gfpga === ejection_channels_112__bench) && !(ejection_channels_112__bench === 1'bx)) begin
				ejection_channels_112__flag <= 1'b1;
			end else begin
				ejection_channels_112__flag<= 1'b0;
			end
			if(!(ejection_channels_111__gfpga === ejection_channels_111__bench) && !(ejection_channels_111__bench === 1'bx)) begin
				ejection_channels_111__flag <= 1'b1;
			end else begin
				ejection_channels_111__flag<= 1'b0;
			end
			if(!(ejection_channels_110__gfpga === ejection_channels_110__bench) && !(ejection_channels_110__bench === 1'bx)) begin
				ejection_channels_110__flag <= 1'b1;
			end else begin
				ejection_channels_110__flag<= 1'b0;
			end
			if(!(ejection_channels_109__gfpga === ejection_channels_109__bench) && !(ejection_channels_109__bench === 1'bx)) begin
				ejection_channels_109__flag <= 1'b1;
			end else begin
				ejection_channels_109__flag<= 1'b0;
			end
			if(!(ejection_channels_108__gfpga === ejection_channels_108__bench) && !(ejection_channels_108__bench === 1'bx)) begin
				ejection_channels_108__flag <= 1'b1;
			end else begin
				ejection_channels_108__flag<= 1'b0;
			end
			if(!(ejection_channels_107__gfpga === ejection_channels_107__bench) && !(ejection_channels_107__bench === 1'bx)) begin
				ejection_channels_107__flag <= 1'b1;
			end else begin
				ejection_channels_107__flag<= 1'b0;
			end
			if(!(ejection_channels_106__gfpga === ejection_channels_106__bench) && !(ejection_channels_106__bench === 1'bx)) begin
				ejection_channels_106__flag <= 1'b1;
			end else begin
				ejection_channels_106__flag<= 1'b0;
			end
			if(!(ejection_channels_105__gfpga === ejection_channels_105__bench) && !(ejection_channels_105__bench === 1'bx)) begin
				ejection_channels_105__flag <= 1'b1;
			end else begin
				ejection_channels_105__flag<= 1'b0;
			end
			if(!(ejection_channels_104__gfpga === ejection_channels_104__bench) && !(ejection_channels_104__bench === 1'bx)) begin
				ejection_channels_104__flag <= 1'b1;
			end else begin
				ejection_channels_104__flag<= 1'b0;
			end
			if(!(ejection_channels_103__gfpga === ejection_channels_103__bench) && !(ejection_channels_103__bench === 1'bx)) begin
				ejection_channels_103__flag <= 1'b1;
			end else begin
				ejection_channels_103__flag<= 1'b0;
			end
			if(!(ejection_channels_102__gfpga === ejection_channels_102__bench) && !(ejection_channels_102__bench === 1'bx)) begin
				ejection_channels_102__flag <= 1'b1;
			end else begin
				ejection_channels_102__flag<= 1'b0;
			end
			if(!(ejection_channels_101__gfpga === ejection_channels_101__bench) && !(ejection_channels_101__bench === 1'bx)) begin
				ejection_channels_101__flag <= 1'b1;
			end else begin
				ejection_channels_101__flag<= 1'b0;
			end
			if(!(ejection_channels_100__gfpga === ejection_channels_100__bench) && !(ejection_channels_100__bench === 1'bx)) begin
				ejection_channels_100__flag <= 1'b1;
			end else begin
				ejection_channels_100__flag<= 1'b0;
			end
			if(!(ejection_channels_99__gfpga === ejection_channels_99__bench) && !(ejection_channels_99__bench === 1'bx)) begin
				ejection_channels_99__flag <= 1'b1;
			end else begin
				ejection_channels_99__flag<= 1'b0;
			end
			if(!(ejection_channels_98__gfpga === ejection_channels_98__bench) && !(ejection_channels_98__bench === 1'bx)) begin
				ejection_channels_98__flag <= 1'b1;
			end else begin
				ejection_channels_98__flag<= 1'b0;
			end
			if(!(ejection_channels_97__gfpga === ejection_channels_97__bench) && !(ejection_channels_97__bench === 1'bx)) begin
				ejection_channels_97__flag <= 1'b1;
			end else begin
				ejection_channels_97__flag<= 1'b0;
			end
			if(!(ejection_channels_96__gfpga === ejection_channels_96__bench) && !(ejection_channels_96__bench === 1'bx)) begin
				ejection_channels_96__flag <= 1'b1;
			end else begin
				ejection_channels_96__flag<= 1'b0;
			end
			if(!(ejection_channels_95__gfpga === ejection_channels_95__bench) && !(ejection_channels_95__bench === 1'bx)) begin
				ejection_channels_95__flag <= 1'b1;
			end else begin
				ejection_channels_95__flag<= 1'b0;
			end
			if(!(ejection_channels_94__gfpga === ejection_channels_94__bench) && !(ejection_channels_94__bench === 1'bx)) begin
				ejection_channels_94__flag <= 1'b1;
			end else begin
				ejection_channels_94__flag<= 1'b0;
			end
			if(!(ejection_channels_93__gfpga === ejection_channels_93__bench) && !(ejection_channels_93__bench === 1'bx)) begin
				ejection_channels_93__flag <= 1'b1;
			end else begin
				ejection_channels_93__flag<= 1'b0;
			end
			if(!(ejection_channels_92__gfpga === ejection_channels_92__bench) && !(ejection_channels_92__bench === 1'bx)) begin
				ejection_channels_92__flag <= 1'b1;
			end else begin
				ejection_channels_92__flag<= 1'b0;
			end
			if(!(ejection_channels_91__gfpga === ejection_channels_91__bench) && !(ejection_channels_91__bench === 1'bx)) begin
				ejection_channels_91__flag <= 1'b1;
			end else begin
				ejection_channels_91__flag<= 1'b0;
			end
			if(!(ejection_channels_90__gfpga === ejection_channels_90__bench) && !(ejection_channels_90__bench === 1'bx)) begin
				ejection_channels_90__flag <= 1'b1;
			end else begin
				ejection_channels_90__flag<= 1'b0;
			end
			if(!(ejection_channels_89__gfpga === ejection_channels_89__bench) && !(ejection_channels_89__bench === 1'bx)) begin
				ejection_channels_89__flag <= 1'b1;
			end else begin
				ejection_channels_89__flag<= 1'b0;
			end
			if(!(ejection_channels_88__gfpga === ejection_channels_88__bench) && !(ejection_channels_88__bench === 1'bx)) begin
				ejection_channels_88__flag <= 1'b1;
			end else begin
				ejection_channels_88__flag<= 1'b0;
			end
			if(!(ejection_channels_87__gfpga === ejection_channels_87__bench) && !(ejection_channels_87__bench === 1'bx)) begin
				ejection_channels_87__flag <= 1'b1;
			end else begin
				ejection_channels_87__flag<= 1'b0;
			end
			if(!(ejection_channels_86__gfpga === ejection_channels_86__bench) && !(ejection_channels_86__bench === 1'bx)) begin
				ejection_channels_86__flag <= 1'b1;
			end else begin
				ejection_channels_86__flag<= 1'b0;
			end
			if(!(ejection_channels_85__gfpga === ejection_channels_85__bench) && !(ejection_channels_85__bench === 1'bx)) begin
				ejection_channels_85__flag <= 1'b1;
			end else begin
				ejection_channels_85__flag<= 1'b0;
			end
			if(!(ejection_channels_84__gfpga === ejection_channels_84__bench) && !(ejection_channels_84__bench === 1'bx)) begin
				ejection_channels_84__flag <= 1'b1;
			end else begin
				ejection_channels_84__flag<= 1'b0;
			end
			if(!(ejection_channels_83__gfpga === ejection_channels_83__bench) && !(ejection_channels_83__bench === 1'bx)) begin
				ejection_channels_83__flag <= 1'b1;
			end else begin
				ejection_channels_83__flag<= 1'b0;
			end
			if(!(ejection_channels_82__gfpga === ejection_channels_82__bench) && !(ejection_channels_82__bench === 1'bx)) begin
				ejection_channels_82__flag <= 1'b1;
			end else begin
				ejection_channels_82__flag<= 1'b0;
			end
			if(!(ejection_channels_81__gfpga === ejection_channels_81__bench) && !(ejection_channels_81__bench === 1'bx)) begin
				ejection_channels_81__flag <= 1'b1;
			end else begin
				ejection_channels_81__flag<= 1'b0;
			end
			if(!(ejection_channels_80__gfpga === ejection_channels_80__bench) && !(ejection_channels_80__bench === 1'bx)) begin
				ejection_channels_80__flag <= 1'b1;
			end else begin
				ejection_channels_80__flag<= 1'b0;
			end
			if(!(ejection_channels_79__gfpga === ejection_channels_79__bench) && !(ejection_channels_79__bench === 1'bx)) begin
				ejection_channels_79__flag <= 1'b1;
			end else begin
				ejection_channels_79__flag<= 1'b0;
			end
			if(!(ejection_channels_78__gfpga === ejection_channels_78__bench) && !(ejection_channels_78__bench === 1'bx)) begin
				ejection_channels_78__flag <= 1'b1;
			end else begin
				ejection_channels_78__flag<= 1'b0;
			end
			if(!(ejection_channels_77__gfpga === ejection_channels_77__bench) && !(ejection_channels_77__bench === 1'bx)) begin
				ejection_channels_77__flag <= 1'b1;
			end else begin
				ejection_channels_77__flag<= 1'b0;
			end
			if(!(ejection_channels_76__gfpga === ejection_channels_76__bench) && !(ejection_channels_76__bench === 1'bx)) begin
				ejection_channels_76__flag <= 1'b1;
			end else begin
				ejection_channels_76__flag<= 1'b0;
			end
			if(!(ejection_channels_75__gfpga === ejection_channels_75__bench) && !(ejection_channels_75__bench === 1'bx)) begin
				ejection_channels_75__flag <= 1'b1;
			end else begin
				ejection_channels_75__flag<= 1'b0;
			end
			if(!(ejection_channels_74__gfpga === ejection_channels_74__bench) && !(ejection_channels_74__bench === 1'bx)) begin
				ejection_channels_74__flag <= 1'b1;
			end else begin
				ejection_channels_74__flag<= 1'b0;
			end
			if(!(ejection_channels_73__gfpga === ejection_channels_73__bench) && !(ejection_channels_73__bench === 1'bx)) begin
				ejection_channels_73__flag <= 1'b1;
			end else begin
				ejection_channels_73__flag<= 1'b0;
			end
			if(!(ejection_channels_72__gfpga === ejection_channels_72__bench) && !(ejection_channels_72__bench === 1'bx)) begin
				ejection_channels_72__flag <= 1'b1;
			end else begin
				ejection_channels_72__flag<= 1'b0;
			end
			if(!(ejection_channels_71__gfpga === ejection_channels_71__bench) && !(ejection_channels_71__bench === 1'bx)) begin
				ejection_channels_71__flag <= 1'b1;
			end else begin
				ejection_channels_71__flag<= 1'b0;
			end
			if(!(ejection_channels_70__gfpga === ejection_channels_70__bench) && !(ejection_channels_70__bench === 1'bx)) begin
				ejection_channels_70__flag <= 1'b1;
			end else begin
				ejection_channels_70__flag<= 1'b0;
			end
			if(!(ejection_channels_69__gfpga === ejection_channels_69__bench) && !(ejection_channels_69__bench === 1'bx)) begin
				ejection_channels_69__flag <= 1'b1;
			end else begin
				ejection_channels_69__flag<= 1'b0;
			end
			if(!(ejection_channels_68__gfpga === ejection_channels_68__bench) && !(ejection_channels_68__bench === 1'bx)) begin
				ejection_channels_68__flag <= 1'b1;
			end else begin
				ejection_channels_68__flag<= 1'b0;
			end
			if(!(ejection_channels_67__gfpga === ejection_channels_67__bench) && !(ejection_channels_67__bench === 1'bx)) begin
				ejection_channels_67__flag <= 1'b1;
			end else begin
				ejection_channels_67__flag<= 1'b0;
			end
			if(!(ejection_channels_66__gfpga === ejection_channels_66__bench) && !(ejection_channels_66__bench === 1'bx)) begin
				ejection_channels_66__flag <= 1'b1;
			end else begin
				ejection_channels_66__flag<= 1'b0;
			end
			if(!(ejection_channels_65__gfpga === ejection_channels_65__bench) && !(ejection_channels_65__bench === 1'bx)) begin
				ejection_channels_65__flag <= 1'b1;
			end else begin
				ejection_channels_65__flag<= 1'b0;
			end
			if(!(ejection_channels_64__gfpga === ejection_channels_64__bench) && !(ejection_channels_64__bench === 1'bx)) begin
				ejection_channels_64__flag <= 1'b1;
			end else begin
				ejection_channels_64__flag<= 1'b0;
			end
			if(!(ejection_channels_63__gfpga === ejection_channels_63__bench) && !(ejection_channels_63__bench === 1'bx)) begin
				ejection_channels_63__flag <= 1'b1;
			end else begin
				ejection_channels_63__flag<= 1'b0;
			end
			if(!(ejection_channels_62__gfpga === ejection_channels_62__bench) && !(ejection_channels_62__bench === 1'bx)) begin
				ejection_channels_62__flag <= 1'b1;
			end else begin
				ejection_channels_62__flag<= 1'b0;
			end
			if(!(ejection_channels_61__gfpga === ejection_channels_61__bench) && !(ejection_channels_61__bench === 1'bx)) begin
				ejection_channels_61__flag <= 1'b1;
			end else begin
				ejection_channels_61__flag<= 1'b0;
			end
			if(!(ejection_channels_60__gfpga === ejection_channels_60__bench) && !(ejection_channels_60__bench === 1'bx)) begin
				ejection_channels_60__flag <= 1'b1;
			end else begin
				ejection_channels_60__flag<= 1'b0;
			end
			if(!(ejection_channels_59__gfpga === ejection_channels_59__bench) && !(ejection_channels_59__bench === 1'bx)) begin
				ejection_channels_59__flag <= 1'b1;
			end else begin
				ejection_channels_59__flag<= 1'b0;
			end
			if(!(ejection_channels_58__gfpga === ejection_channels_58__bench) && !(ejection_channels_58__bench === 1'bx)) begin
				ejection_channels_58__flag <= 1'b1;
			end else begin
				ejection_channels_58__flag<= 1'b0;
			end
			if(!(ejection_channels_57__gfpga === ejection_channels_57__bench) && !(ejection_channels_57__bench === 1'bx)) begin
				ejection_channels_57__flag <= 1'b1;
			end else begin
				ejection_channels_57__flag<= 1'b0;
			end
			if(!(ejection_channels_56__gfpga === ejection_channels_56__bench) && !(ejection_channels_56__bench === 1'bx)) begin
				ejection_channels_56__flag <= 1'b1;
			end else begin
				ejection_channels_56__flag<= 1'b0;
			end
			if(!(ejection_channels_55__gfpga === ejection_channels_55__bench) && !(ejection_channels_55__bench === 1'bx)) begin
				ejection_channels_55__flag <= 1'b1;
			end else begin
				ejection_channels_55__flag<= 1'b0;
			end
			if(!(ejection_channels_54__gfpga === ejection_channels_54__bench) && !(ejection_channels_54__bench === 1'bx)) begin
				ejection_channels_54__flag <= 1'b1;
			end else begin
				ejection_channels_54__flag<= 1'b0;
			end
			if(!(ejection_channels_53__gfpga === ejection_channels_53__bench) && !(ejection_channels_53__bench === 1'bx)) begin
				ejection_channels_53__flag <= 1'b1;
			end else begin
				ejection_channels_53__flag<= 1'b0;
			end
			if(!(ejection_channels_52__gfpga === ejection_channels_52__bench) && !(ejection_channels_52__bench === 1'bx)) begin
				ejection_channels_52__flag <= 1'b1;
			end else begin
				ejection_channels_52__flag<= 1'b0;
			end
			if(!(ejection_channels_51__gfpga === ejection_channels_51__bench) && !(ejection_channels_51__bench === 1'bx)) begin
				ejection_channels_51__flag <= 1'b1;
			end else begin
				ejection_channels_51__flag<= 1'b0;
			end
			if(!(ejection_channels_50__gfpga === ejection_channels_50__bench) && !(ejection_channels_50__bench === 1'bx)) begin
				ejection_channels_50__flag <= 1'b1;
			end else begin
				ejection_channels_50__flag<= 1'b0;
			end
			if(!(ejection_channels_49__gfpga === ejection_channels_49__bench) && !(ejection_channels_49__bench === 1'bx)) begin
				ejection_channels_49__flag <= 1'b1;
			end else begin
				ejection_channels_49__flag<= 1'b0;
			end
			if(!(ejection_channels_48__gfpga === ejection_channels_48__bench) && !(ejection_channels_48__bench === 1'bx)) begin
				ejection_channels_48__flag <= 1'b1;
			end else begin
				ejection_channels_48__flag<= 1'b0;
			end
			if(!(ejection_channels_47__gfpga === ejection_channels_47__bench) && !(ejection_channels_47__bench === 1'bx)) begin
				ejection_channels_47__flag <= 1'b1;
			end else begin
				ejection_channels_47__flag<= 1'b0;
			end
			if(!(ejection_channels_46__gfpga === ejection_channels_46__bench) && !(ejection_channels_46__bench === 1'bx)) begin
				ejection_channels_46__flag <= 1'b1;
			end else begin
				ejection_channels_46__flag<= 1'b0;
			end
			if(!(ejection_channels_45__gfpga === ejection_channels_45__bench) && !(ejection_channels_45__bench === 1'bx)) begin
				ejection_channels_45__flag <= 1'b1;
			end else begin
				ejection_channels_45__flag<= 1'b0;
			end
			if(!(ejection_channels_44__gfpga === ejection_channels_44__bench) && !(ejection_channels_44__bench === 1'bx)) begin
				ejection_channels_44__flag <= 1'b1;
			end else begin
				ejection_channels_44__flag<= 1'b0;
			end
			if(!(ejection_channels_43__gfpga === ejection_channels_43__bench) && !(ejection_channels_43__bench === 1'bx)) begin
				ejection_channels_43__flag <= 1'b1;
			end else begin
				ejection_channels_43__flag<= 1'b0;
			end
			if(!(ejection_channels_42__gfpga === ejection_channels_42__bench) && !(ejection_channels_42__bench === 1'bx)) begin
				ejection_channels_42__flag <= 1'b1;
			end else begin
				ejection_channels_42__flag<= 1'b0;
			end
			if(!(ejection_channels_41__gfpga === ejection_channels_41__bench) && !(ejection_channels_41__bench === 1'bx)) begin
				ejection_channels_41__flag <= 1'b1;
			end else begin
				ejection_channels_41__flag<= 1'b0;
			end
			if(!(ejection_channels_40__gfpga === ejection_channels_40__bench) && !(ejection_channels_40__bench === 1'bx)) begin
				ejection_channels_40__flag <= 1'b1;
			end else begin
				ejection_channels_40__flag<= 1'b0;
			end
			if(!(ejection_channels_39__gfpga === ejection_channels_39__bench) && !(ejection_channels_39__bench === 1'bx)) begin
				ejection_channels_39__flag <= 1'b1;
			end else begin
				ejection_channels_39__flag<= 1'b0;
			end
			if(!(ejection_channels_38__gfpga === ejection_channels_38__bench) && !(ejection_channels_38__bench === 1'bx)) begin
				ejection_channels_38__flag <= 1'b1;
			end else begin
				ejection_channels_38__flag<= 1'b0;
			end
			if(!(ejection_channels_37__gfpga === ejection_channels_37__bench) && !(ejection_channels_37__bench === 1'bx)) begin
				ejection_channels_37__flag <= 1'b1;
			end else begin
				ejection_channels_37__flag<= 1'b0;
			end
			if(!(ejection_channels_36__gfpga === ejection_channels_36__bench) && !(ejection_channels_36__bench === 1'bx)) begin
				ejection_channels_36__flag <= 1'b1;
			end else begin
				ejection_channels_36__flag<= 1'b0;
			end
			if(!(ejection_channels_35__gfpga === ejection_channels_35__bench) && !(ejection_channels_35__bench === 1'bx)) begin
				ejection_channels_35__flag <= 1'b1;
			end else begin
				ejection_channels_35__flag<= 1'b0;
			end
			if(!(ejection_channels_34__gfpga === ejection_channels_34__bench) && !(ejection_channels_34__bench === 1'bx)) begin
				ejection_channels_34__flag <= 1'b1;
			end else begin
				ejection_channels_34__flag<= 1'b0;
			end
			if(!(ejection_channels_33__gfpga === ejection_channels_33__bench) && !(ejection_channels_33__bench === 1'bx)) begin
				ejection_channels_33__flag <= 1'b1;
			end else begin
				ejection_channels_33__flag<= 1'b0;
			end
			if(!(ejection_channels_32__gfpga === ejection_channels_32__bench) && !(ejection_channels_32__bench === 1'bx)) begin
				ejection_channels_32__flag <= 1'b1;
			end else begin
				ejection_channels_32__flag<= 1'b0;
			end
			if(!(ejection_channels_31__gfpga === ejection_channels_31__bench) && !(ejection_channels_31__bench === 1'bx)) begin
				ejection_channels_31__flag <= 1'b1;
			end else begin
				ejection_channels_31__flag<= 1'b0;
			end
			if(!(ejection_channels_30__gfpga === ejection_channels_30__bench) && !(ejection_channels_30__bench === 1'bx)) begin
				ejection_channels_30__flag <= 1'b1;
			end else begin
				ejection_channels_30__flag<= 1'b0;
			end
			if(!(ejection_channels_29__gfpga === ejection_channels_29__bench) && !(ejection_channels_29__bench === 1'bx)) begin
				ejection_channels_29__flag <= 1'b1;
			end else begin
				ejection_channels_29__flag<= 1'b0;
			end
			if(!(ejection_channels_28__gfpga === ejection_channels_28__bench) && !(ejection_channels_28__bench === 1'bx)) begin
				ejection_channels_28__flag <= 1'b1;
			end else begin
				ejection_channels_28__flag<= 1'b0;
			end
			if(!(ejection_channels_27__gfpga === ejection_channels_27__bench) && !(ejection_channels_27__bench === 1'bx)) begin
				ejection_channels_27__flag <= 1'b1;
			end else begin
				ejection_channels_27__flag<= 1'b0;
			end
			if(!(ejection_channels_26__gfpga === ejection_channels_26__bench) && !(ejection_channels_26__bench === 1'bx)) begin
				ejection_channels_26__flag <= 1'b1;
			end else begin
				ejection_channels_26__flag<= 1'b0;
			end
			if(!(ejection_channels_25__gfpga === ejection_channels_25__bench) && !(ejection_channels_25__bench === 1'bx)) begin
				ejection_channels_25__flag <= 1'b1;
			end else begin
				ejection_channels_25__flag<= 1'b0;
			end
			if(!(ejection_channels_24__gfpga === ejection_channels_24__bench) && !(ejection_channels_24__bench === 1'bx)) begin
				ejection_channels_24__flag <= 1'b1;
			end else begin
				ejection_channels_24__flag<= 1'b0;
			end
			if(!(ejection_channels_23__gfpga === ejection_channels_23__bench) && !(ejection_channels_23__bench === 1'bx)) begin
				ejection_channels_23__flag <= 1'b1;
			end else begin
				ejection_channels_23__flag<= 1'b0;
			end
			if(!(ejection_channels_22__gfpga === ejection_channels_22__bench) && !(ejection_channels_22__bench === 1'bx)) begin
				ejection_channels_22__flag <= 1'b1;
			end else begin
				ejection_channels_22__flag<= 1'b0;
			end
			if(!(ejection_channels_21__gfpga === ejection_channels_21__bench) && !(ejection_channels_21__bench === 1'bx)) begin
				ejection_channels_21__flag <= 1'b1;
			end else begin
				ejection_channels_21__flag<= 1'b0;
			end
			if(!(ejection_channels_20__gfpga === ejection_channels_20__bench) && !(ejection_channels_20__bench === 1'bx)) begin
				ejection_channels_20__flag <= 1'b1;
			end else begin
				ejection_channels_20__flag<= 1'b0;
			end
			if(!(ejection_channels_19__gfpga === ejection_channels_19__bench) && !(ejection_channels_19__bench === 1'bx)) begin
				ejection_channels_19__flag <= 1'b1;
			end else begin
				ejection_channels_19__flag<= 1'b0;
			end
			if(!(ejection_channels_18__gfpga === ejection_channels_18__bench) && !(ejection_channels_18__bench === 1'bx)) begin
				ejection_channels_18__flag <= 1'b1;
			end else begin
				ejection_channels_18__flag<= 1'b0;
			end
			if(!(ejection_channels_17__gfpga === ejection_channels_17__bench) && !(ejection_channels_17__bench === 1'bx)) begin
				ejection_channels_17__flag <= 1'b1;
			end else begin
				ejection_channels_17__flag<= 1'b0;
			end
			if(!(ejection_channels_16__gfpga === ejection_channels_16__bench) && !(ejection_channels_16__bench === 1'bx)) begin
				ejection_channels_16__flag <= 1'b1;
			end else begin
				ejection_channels_16__flag<= 1'b0;
			end
			if(!(ejection_channels_15__gfpga === ejection_channels_15__bench) && !(ejection_channels_15__bench === 1'bx)) begin
				ejection_channels_15__flag <= 1'b1;
			end else begin
				ejection_channels_15__flag<= 1'b0;
			end
			if(!(ejection_channels_14__gfpga === ejection_channels_14__bench) && !(ejection_channels_14__bench === 1'bx)) begin
				ejection_channels_14__flag <= 1'b1;
			end else begin
				ejection_channels_14__flag<= 1'b0;
			end
			if(!(ejection_channels_13__gfpga === ejection_channels_13__bench) && !(ejection_channels_13__bench === 1'bx)) begin
				ejection_channels_13__flag <= 1'b1;
			end else begin
				ejection_channels_13__flag<= 1'b0;
			end
			if(!(ejection_channels_12__gfpga === ejection_channels_12__bench) && !(ejection_channels_12__bench === 1'bx)) begin
				ejection_channels_12__flag <= 1'b1;
			end else begin
				ejection_channels_12__flag<= 1'b0;
			end
			if(!(ejection_channels_11__gfpga === ejection_channels_11__bench) && !(ejection_channels_11__bench === 1'bx)) begin
				ejection_channels_11__flag <= 1'b1;
			end else begin
				ejection_channels_11__flag<= 1'b0;
			end
			if(!(ejection_channels_10__gfpga === ejection_channels_10__bench) && !(ejection_channels_10__bench === 1'bx)) begin
				ejection_channels_10__flag <= 1'b1;
			end else begin
				ejection_channels_10__flag<= 1'b0;
			end
			if(!(ejection_channels_9__gfpga === ejection_channels_9__bench) && !(ejection_channels_9__bench === 1'bx)) begin
				ejection_channels_9__flag <= 1'b1;
			end else begin
				ejection_channels_9__flag<= 1'b0;
			end
			if(!(ejection_channels_8__gfpga === ejection_channels_8__bench) && !(ejection_channels_8__bench === 1'bx)) begin
				ejection_channels_8__flag <= 1'b1;
			end else begin
				ejection_channels_8__flag<= 1'b0;
			end
			if(!(ejection_channels_7__gfpga === ejection_channels_7__bench) && !(ejection_channels_7__bench === 1'bx)) begin
				ejection_channels_7__flag <= 1'b1;
			end else begin
				ejection_channels_7__flag<= 1'b0;
			end
			if(!(ejection_channels_6__gfpga === ejection_channels_6__bench) && !(ejection_channels_6__bench === 1'bx)) begin
				ejection_channels_6__flag <= 1'b1;
			end else begin
				ejection_channels_6__flag<= 1'b0;
			end
			if(!(ejection_channels_5__gfpga === ejection_channels_5__bench) && !(ejection_channels_5__bench === 1'bx)) begin
				ejection_channels_5__flag <= 1'b1;
			end else begin
				ejection_channels_5__flag<= 1'b0;
			end
			if(!(ejection_channels_4__gfpga === ejection_channels_4__bench) && !(ejection_channels_4__bench === 1'bx)) begin
				ejection_channels_4__flag <= 1'b1;
			end else begin
				ejection_channels_4__flag<= 1'b0;
			end
			if(!(ejection_channels_3__gfpga === ejection_channels_3__bench) && !(ejection_channels_3__bench === 1'bx)) begin
				ejection_channels_3__flag <= 1'b1;
			end else begin
				ejection_channels_3__flag<= 1'b0;
			end
			if(!(ejection_channels_2__gfpga === ejection_channels_2__bench) && !(ejection_channels_2__bench === 1'bx)) begin
				ejection_channels_2__flag <= 1'b1;
			end else begin
				ejection_channels_2__flag<= 1'b0;
			end
			if(!(ejection_channels_1__gfpga === ejection_channels_1__bench) && !(ejection_channels_1__bench === 1'bx)) begin
				ejection_channels_1__flag <= 1'b1;
			end else begin
				ejection_channels_1__flag<= 1'b0;
			end
			if(!(ejection_channels_0__gfpga === ejection_channels_0__bench) && !(ejection_channels_0__bench === 1'bx)) begin
				ejection_channels_0__flag <= 1'b1;
			end else begin
				ejection_channels_0__flag<= 1'b0;
			end
			if(!(rtr_error_8__gfpga === rtr_error_8__bench) && !(rtr_error_8__bench === 1'bx)) begin
				rtr_error_8__flag <= 1'b1;
			end else begin
				rtr_error_8__flag<= 1'b0;
			end
			if(!(rtr_error_7__gfpga === rtr_error_7__bench) && !(rtr_error_7__bench === 1'bx)) begin
				rtr_error_7__flag <= 1'b1;
			end else begin
				rtr_error_7__flag<= 1'b0;
			end
			if(!(rtr_error_6__gfpga === rtr_error_6__bench) && !(rtr_error_6__bench === 1'bx)) begin
				rtr_error_6__flag <= 1'b1;
			end else begin
				rtr_error_6__flag<= 1'b0;
			end
			if(!(rtr_error_5__gfpga === rtr_error_5__bench) && !(rtr_error_5__bench === 1'bx)) begin
				rtr_error_5__flag <= 1'b1;
			end else begin
				rtr_error_5__flag<= 1'b0;
			end
			if(!(rtr_error_4__gfpga === rtr_error_4__bench) && !(rtr_error_4__bench === 1'bx)) begin
				rtr_error_4__flag <= 1'b1;
			end else begin
				rtr_error_4__flag<= 1'b0;
			end
			if(!(rtr_error_3__gfpga === rtr_error_3__bench) && !(rtr_error_3__bench === 1'bx)) begin
				rtr_error_3__flag <= 1'b1;
			end else begin
				rtr_error_3__flag<= 1'b0;
			end
			if(!(rtr_error_2__gfpga === rtr_error_2__bench) && !(rtr_error_2__bench === 1'bx)) begin
				rtr_error_2__flag <= 1'b1;
			end else begin
				rtr_error_2__flag<= 1'b0;
			end
			if(!(rtr_error_1__gfpga === rtr_error_1__bench) && !(rtr_error_1__bench === 1'bx)) begin
				rtr_error_1__flag <= 1'b1;
			end else begin
				rtr_error_1__flag<= 1'b0;
			end
			if(!(rtr_error_0__gfpga === rtr_error_0__bench) && !(rtr_error_0__bench === 1'bx)) begin
				rtr_error_0__flag <= 1'b1;
			end else begin
				rtr_error_0__flag<= 1'b0;
			end
		end
	end

	always@(posedge injection_flow_ctrl_26__flag) begin
		if(injection_flow_ctrl_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_25__flag) begin
		if(injection_flow_ctrl_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_24__flag) begin
		if(injection_flow_ctrl_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_23__flag) begin
		if(injection_flow_ctrl_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_22__flag) begin
		if(injection_flow_ctrl_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_21__flag) begin
		if(injection_flow_ctrl_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_20__flag) begin
		if(injection_flow_ctrl_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_19__flag) begin
		if(injection_flow_ctrl_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_18__flag) begin
		if(injection_flow_ctrl_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_17__flag) begin
		if(injection_flow_ctrl_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_16__flag) begin
		if(injection_flow_ctrl_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_15__flag) begin
		if(injection_flow_ctrl_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_14__flag) begin
		if(injection_flow_ctrl_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_13__flag) begin
		if(injection_flow_ctrl_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_12__flag) begin
		if(injection_flow_ctrl_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_11__flag) begin
		if(injection_flow_ctrl_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_10__flag) begin
		if(injection_flow_ctrl_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_9__flag) begin
		if(injection_flow_ctrl_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_8__flag) begin
		if(injection_flow_ctrl_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_7__flag) begin
		if(injection_flow_ctrl_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_6__flag) begin
		if(injection_flow_ctrl_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_5__flag) begin
		if(injection_flow_ctrl_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_4__flag) begin
		if(injection_flow_ctrl_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_3__flag) begin
		if(injection_flow_ctrl_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_2__flag) begin
		if(injection_flow_ctrl_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_1__flag) begin
		if(injection_flow_ctrl_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge injection_flow_ctrl_0__flag) begin
		if(injection_flow_ctrl_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on injection_flow_ctrl_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_629__flag) begin
		if(ejection_channels_629__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_629__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_628__flag) begin
		if(ejection_channels_628__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_628__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_627__flag) begin
		if(ejection_channels_627__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_627__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_626__flag) begin
		if(ejection_channels_626__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_626__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_625__flag) begin
		if(ejection_channels_625__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_625__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_624__flag) begin
		if(ejection_channels_624__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_624__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_623__flag) begin
		if(ejection_channels_623__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_623__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_622__flag) begin
		if(ejection_channels_622__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_622__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_621__flag) begin
		if(ejection_channels_621__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_621__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_620__flag) begin
		if(ejection_channels_620__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_620__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_619__flag) begin
		if(ejection_channels_619__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_619__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_618__flag) begin
		if(ejection_channels_618__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_618__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_617__flag) begin
		if(ejection_channels_617__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_617__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_616__flag) begin
		if(ejection_channels_616__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_616__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_615__flag) begin
		if(ejection_channels_615__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_615__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_614__flag) begin
		if(ejection_channels_614__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_614__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_613__flag) begin
		if(ejection_channels_613__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_613__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_612__flag) begin
		if(ejection_channels_612__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_612__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_611__flag) begin
		if(ejection_channels_611__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_611__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_610__flag) begin
		if(ejection_channels_610__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_610__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_609__flag) begin
		if(ejection_channels_609__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_609__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_608__flag) begin
		if(ejection_channels_608__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_608__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_607__flag) begin
		if(ejection_channels_607__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_607__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_606__flag) begin
		if(ejection_channels_606__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_606__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_605__flag) begin
		if(ejection_channels_605__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_605__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_604__flag) begin
		if(ejection_channels_604__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_604__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_603__flag) begin
		if(ejection_channels_603__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_603__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_602__flag) begin
		if(ejection_channels_602__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_602__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_601__flag) begin
		if(ejection_channels_601__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_601__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_600__flag) begin
		if(ejection_channels_600__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_600__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_599__flag) begin
		if(ejection_channels_599__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_599__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_598__flag) begin
		if(ejection_channels_598__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_598__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_597__flag) begin
		if(ejection_channels_597__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_597__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_596__flag) begin
		if(ejection_channels_596__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_596__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_595__flag) begin
		if(ejection_channels_595__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_595__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_594__flag) begin
		if(ejection_channels_594__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_594__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_593__flag) begin
		if(ejection_channels_593__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_593__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_592__flag) begin
		if(ejection_channels_592__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_592__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_591__flag) begin
		if(ejection_channels_591__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_591__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_590__flag) begin
		if(ejection_channels_590__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_590__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_589__flag) begin
		if(ejection_channels_589__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_589__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_588__flag) begin
		if(ejection_channels_588__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_588__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_587__flag) begin
		if(ejection_channels_587__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_587__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_586__flag) begin
		if(ejection_channels_586__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_586__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_585__flag) begin
		if(ejection_channels_585__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_585__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_584__flag) begin
		if(ejection_channels_584__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_584__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_583__flag) begin
		if(ejection_channels_583__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_583__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_582__flag) begin
		if(ejection_channels_582__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_582__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_581__flag) begin
		if(ejection_channels_581__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_581__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_580__flag) begin
		if(ejection_channels_580__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_580__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_579__flag) begin
		if(ejection_channels_579__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_579__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_578__flag) begin
		if(ejection_channels_578__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_578__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_577__flag) begin
		if(ejection_channels_577__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_577__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_576__flag) begin
		if(ejection_channels_576__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_576__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_575__flag) begin
		if(ejection_channels_575__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_575__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_574__flag) begin
		if(ejection_channels_574__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_574__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_573__flag) begin
		if(ejection_channels_573__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_573__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_572__flag) begin
		if(ejection_channels_572__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_572__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_571__flag) begin
		if(ejection_channels_571__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_571__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_570__flag) begin
		if(ejection_channels_570__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_570__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_569__flag) begin
		if(ejection_channels_569__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_569__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_568__flag) begin
		if(ejection_channels_568__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_568__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_567__flag) begin
		if(ejection_channels_567__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_567__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_566__flag) begin
		if(ejection_channels_566__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_566__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_565__flag) begin
		if(ejection_channels_565__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_565__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_564__flag) begin
		if(ejection_channels_564__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_564__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_563__flag) begin
		if(ejection_channels_563__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_563__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_562__flag) begin
		if(ejection_channels_562__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_562__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_561__flag) begin
		if(ejection_channels_561__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_561__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_560__flag) begin
		if(ejection_channels_560__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_560__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_559__flag) begin
		if(ejection_channels_559__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_559__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_558__flag) begin
		if(ejection_channels_558__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_558__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_557__flag) begin
		if(ejection_channels_557__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_557__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_556__flag) begin
		if(ejection_channels_556__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_556__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_555__flag) begin
		if(ejection_channels_555__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_555__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_554__flag) begin
		if(ejection_channels_554__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_554__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_553__flag) begin
		if(ejection_channels_553__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_553__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_552__flag) begin
		if(ejection_channels_552__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_552__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_551__flag) begin
		if(ejection_channels_551__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_551__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_550__flag) begin
		if(ejection_channels_550__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_550__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_549__flag) begin
		if(ejection_channels_549__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_549__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_548__flag) begin
		if(ejection_channels_548__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_548__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_547__flag) begin
		if(ejection_channels_547__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_547__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_546__flag) begin
		if(ejection_channels_546__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_546__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_545__flag) begin
		if(ejection_channels_545__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_545__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_544__flag) begin
		if(ejection_channels_544__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_544__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_543__flag) begin
		if(ejection_channels_543__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_543__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_542__flag) begin
		if(ejection_channels_542__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_542__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_541__flag) begin
		if(ejection_channels_541__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_541__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_540__flag) begin
		if(ejection_channels_540__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_540__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_539__flag) begin
		if(ejection_channels_539__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_539__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_538__flag) begin
		if(ejection_channels_538__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_538__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_537__flag) begin
		if(ejection_channels_537__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_537__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_536__flag) begin
		if(ejection_channels_536__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_536__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_535__flag) begin
		if(ejection_channels_535__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_535__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_534__flag) begin
		if(ejection_channels_534__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_534__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_533__flag) begin
		if(ejection_channels_533__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_533__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_532__flag) begin
		if(ejection_channels_532__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_532__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_531__flag) begin
		if(ejection_channels_531__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_531__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_530__flag) begin
		if(ejection_channels_530__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_530__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_529__flag) begin
		if(ejection_channels_529__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_529__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_528__flag) begin
		if(ejection_channels_528__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_528__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_527__flag) begin
		if(ejection_channels_527__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_527__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_526__flag) begin
		if(ejection_channels_526__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_526__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_525__flag) begin
		if(ejection_channels_525__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_525__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_524__flag) begin
		if(ejection_channels_524__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_524__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_523__flag) begin
		if(ejection_channels_523__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_523__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_522__flag) begin
		if(ejection_channels_522__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_522__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_521__flag) begin
		if(ejection_channels_521__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_521__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_520__flag) begin
		if(ejection_channels_520__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_520__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_519__flag) begin
		if(ejection_channels_519__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_519__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_518__flag) begin
		if(ejection_channels_518__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_518__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_517__flag) begin
		if(ejection_channels_517__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_517__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_516__flag) begin
		if(ejection_channels_516__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_516__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_515__flag) begin
		if(ejection_channels_515__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_515__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_514__flag) begin
		if(ejection_channels_514__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_514__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_513__flag) begin
		if(ejection_channels_513__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_513__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_512__flag) begin
		if(ejection_channels_512__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_512__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_511__flag) begin
		if(ejection_channels_511__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_511__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_510__flag) begin
		if(ejection_channels_510__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_510__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_509__flag) begin
		if(ejection_channels_509__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_509__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_508__flag) begin
		if(ejection_channels_508__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_508__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_507__flag) begin
		if(ejection_channels_507__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_507__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_506__flag) begin
		if(ejection_channels_506__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_506__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_505__flag) begin
		if(ejection_channels_505__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_505__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_504__flag) begin
		if(ejection_channels_504__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_504__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_503__flag) begin
		if(ejection_channels_503__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_503__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_502__flag) begin
		if(ejection_channels_502__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_502__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_501__flag) begin
		if(ejection_channels_501__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_501__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_500__flag) begin
		if(ejection_channels_500__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_500__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_499__flag) begin
		if(ejection_channels_499__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_499__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_498__flag) begin
		if(ejection_channels_498__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_498__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_497__flag) begin
		if(ejection_channels_497__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_497__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_496__flag) begin
		if(ejection_channels_496__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_496__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_495__flag) begin
		if(ejection_channels_495__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_495__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_494__flag) begin
		if(ejection_channels_494__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_494__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_493__flag) begin
		if(ejection_channels_493__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_493__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_492__flag) begin
		if(ejection_channels_492__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_492__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_491__flag) begin
		if(ejection_channels_491__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_491__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_490__flag) begin
		if(ejection_channels_490__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_490__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_489__flag) begin
		if(ejection_channels_489__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_489__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_488__flag) begin
		if(ejection_channels_488__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_488__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_487__flag) begin
		if(ejection_channels_487__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_487__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_486__flag) begin
		if(ejection_channels_486__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_486__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_485__flag) begin
		if(ejection_channels_485__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_485__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_484__flag) begin
		if(ejection_channels_484__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_484__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_483__flag) begin
		if(ejection_channels_483__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_483__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_482__flag) begin
		if(ejection_channels_482__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_482__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_481__flag) begin
		if(ejection_channels_481__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_481__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_480__flag) begin
		if(ejection_channels_480__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_480__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_479__flag) begin
		if(ejection_channels_479__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_479__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_478__flag) begin
		if(ejection_channels_478__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_478__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_477__flag) begin
		if(ejection_channels_477__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_477__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_476__flag) begin
		if(ejection_channels_476__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_476__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_475__flag) begin
		if(ejection_channels_475__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_475__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_474__flag) begin
		if(ejection_channels_474__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_474__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_473__flag) begin
		if(ejection_channels_473__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_473__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_472__flag) begin
		if(ejection_channels_472__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_472__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_471__flag) begin
		if(ejection_channels_471__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_471__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_470__flag) begin
		if(ejection_channels_470__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_470__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_469__flag) begin
		if(ejection_channels_469__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_469__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_468__flag) begin
		if(ejection_channels_468__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_468__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_467__flag) begin
		if(ejection_channels_467__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_467__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_466__flag) begin
		if(ejection_channels_466__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_466__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_465__flag) begin
		if(ejection_channels_465__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_465__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_464__flag) begin
		if(ejection_channels_464__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_464__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_463__flag) begin
		if(ejection_channels_463__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_463__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_462__flag) begin
		if(ejection_channels_462__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_462__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_461__flag) begin
		if(ejection_channels_461__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_461__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_460__flag) begin
		if(ejection_channels_460__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_460__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_459__flag) begin
		if(ejection_channels_459__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_459__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_458__flag) begin
		if(ejection_channels_458__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_458__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_457__flag) begin
		if(ejection_channels_457__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_457__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_456__flag) begin
		if(ejection_channels_456__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_456__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_455__flag) begin
		if(ejection_channels_455__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_455__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_454__flag) begin
		if(ejection_channels_454__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_454__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_453__flag) begin
		if(ejection_channels_453__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_453__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_452__flag) begin
		if(ejection_channels_452__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_452__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_451__flag) begin
		if(ejection_channels_451__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_451__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_450__flag) begin
		if(ejection_channels_450__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_450__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_449__flag) begin
		if(ejection_channels_449__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_449__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_448__flag) begin
		if(ejection_channels_448__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_448__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_447__flag) begin
		if(ejection_channels_447__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_447__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_446__flag) begin
		if(ejection_channels_446__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_446__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_445__flag) begin
		if(ejection_channels_445__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_445__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_444__flag) begin
		if(ejection_channels_444__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_444__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_443__flag) begin
		if(ejection_channels_443__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_443__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_442__flag) begin
		if(ejection_channels_442__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_442__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_441__flag) begin
		if(ejection_channels_441__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_441__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_440__flag) begin
		if(ejection_channels_440__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_440__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_439__flag) begin
		if(ejection_channels_439__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_439__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_438__flag) begin
		if(ejection_channels_438__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_438__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_437__flag) begin
		if(ejection_channels_437__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_437__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_436__flag) begin
		if(ejection_channels_436__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_436__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_435__flag) begin
		if(ejection_channels_435__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_435__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_434__flag) begin
		if(ejection_channels_434__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_434__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_433__flag) begin
		if(ejection_channels_433__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_433__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_432__flag) begin
		if(ejection_channels_432__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_432__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_431__flag) begin
		if(ejection_channels_431__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_431__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_430__flag) begin
		if(ejection_channels_430__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_430__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_429__flag) begin
		if(ejection_channels_429__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_429__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_428__flag) begin
		if(ejection_channels_428__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_428__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_427__flag) begin
		if(ejection_channels_427__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_427__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_426__flag) begin
		if(ejection_channels_426__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_426__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_425__flag) begin
		if(ejection_channels_425__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_425__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_424__flag) begin
		if(ejection_channels_424__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_424__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_423__flag) begin
		if(ejection_channels_423__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_423__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_422__flag) begin
		if(ejection_channels_422__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_422__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_421__flag) begin
		if(ejection_channels_421__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_421__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_420__flag) begin
		if(ejection_channels_420__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_420__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_419__flag) begin
		if(ejection_channels_419__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_419__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_418__flag) begin
		if(ejection_channels_418__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_418__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_417__flag) begin
		if(ejection_channels_417__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_417__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_416__flag) begin
		if(ejection_channels_416__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_416__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_415__flag) begin
		if(ejection_channels_415__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_415__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_414__flag) begin
		if(ejection_channels_414__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_414__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_413__flag) begin
		if(ejection_channels_413__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_413__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_412__flag) begin
		if(ejection_channels_412__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_412__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_411__flag) begin
		if(ejection_channels_411__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_411__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_410__flag) begin
		if(ejection_channels_410__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_410__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_409__flag) begin
		if(ejection_channels_409__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_409__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_408__flag) begin
		if(ejection_channels_408__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_408__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_407__flag) begin
		if(ejection_channels_407__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_407__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_406__flag) begin
		if(ejection_channels_406__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_406__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_405__flag) begin
		if(ejection_channels_405__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_405__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_404__flag) begin
		if(ejection_channels_404__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_404__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_403__flag) begin
		if(ejection_channels_403__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_403__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_402__flag) begin
		if(ejection_channels_402__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_402__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_401__flag) begin
		if(ejection_channels_401__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_401__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_400__flag) begin
		if(ejection_channels_400__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_400__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_399__flag) begin
		if(ejection_channels_399__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_399__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_398__flag) begin
		if(ejection_channels_398__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_398__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_397__flag) begin
		if(ejection_channels_397__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_397__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_396__flag) begin
		if(ejection_channels_396__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_396__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_395__flag) begin
		if(ejection_channels_395__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_395__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_394__flag) begin
		if(ejection_channels_394__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_394__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_393__flag) begin
		if(ejection_channels_393__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_393__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_392__flag) begin
		if(ejection_channels_392__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_392__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_391__flag) begin
		if(ejection_channels_391__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_391__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_390__flag) begin
		if(ejection_channels_390__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_390__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_389__flag) begin
		if(ejection_channels_389__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_389__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_388__flag) begin
		if(ejection_channels_388__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_388__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_387__flag) begin
		if(ejection_channels_387__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_387__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_386__flag) begin
		if(ejection_channels_386__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_386__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_385__flag) begin
		if(ejection_channels_385__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_385__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_384__flag) begin
		if(ejection_channels_384__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_384__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_383__flag) begin
		if(ejection_channels_383__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_383__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_382__flag) begin
		if(ejection_channels_382__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_382__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_381__flag) begin
		if(ejection_channels_381__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_381__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_380__flag) begin
		if(ejection_channels_380__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_380__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_379__flag) begin
		if(ejection_channels_379__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_379__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_378__flag) begin
		if(ejection_channels_378__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_378__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_377__flag) begin
		if(ejection_channels_377__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_377__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_376__flag) begin
		if(ejection_channels_376__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_376__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_375__flag) begin
		if(ejection_channels_375__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_375__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_374__flag) begin
		if(ejection_channels_374__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_374__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_373__flag) begin
		if(ejection_channels_373__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_373__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_372__flag) begin
		if(ejection_channels_372__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_372__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_371__flag) begin
		if(ejection_channels_371__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_371__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_370__flag) begin
		if(ejection_channels_370__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_370__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_369__flag) begin
		if(ejection_channels_369__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_369__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_368__flag) begin
		if(ejection_channels_368__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_368__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_367__flag) begin
		if(ejection_channels_367__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_367__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_366__flag) begin
		if(ejection_channels_366__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_366__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_365__flag) begin
		if(ejection_channels_365__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_365__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_364__flag) begin
		if(ejection_channels_364__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_364__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_363__flag) begin
		if(ejection_channels_363__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_363__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_362__flag) begin
		if(ejection_channels_362__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_362__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_361__flag) begin
		if(ejection_channels_361__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_361__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_360__flag) begin
		if(ejection_channels_360__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_360__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_359__flag) begin
		if(ejection_channels_359__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_359__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_358__flag) begin
		if(ejection_channels_358__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_358__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_357__flag) begin
		if(ejection_channels_357__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_357__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_356__flag) begin
		if(ejection_channels_356__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_356__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_355__flag) begin
		if(ejection_channels_355__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_355__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_354__flag) begin
		if(ejection_channels_354__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_354__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_353__flag) begin
		if(ejection_channels_353__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_353__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_352__flag) begin
		if(ejection_channels_352__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_352__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_351__flag) begin
		if(ejection_channels_351__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_351__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_350__flag) begin
		if(ejection_channels_350__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_350__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_349__flag) begin
		if(ejection_channels_349__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_349__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_348__flag) begin
		if(ejection_channels_348__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_348__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_347__flag) begin
		if(ejection_channels_347__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_347__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_346__flag) begin
		if(ejection_channels_346__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_346__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_345__flag) begin
		if(ejection_channels_345__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_345__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_344__flag) begin
		if(ejection_channels_344__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_344__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_343__flag) begin
		if(ejection_channels_343__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_343__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_342__flag) begin
		if(ejection_channels_342__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_342__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_341__flag) begin
		if(ejection_channels_341__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_341__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_340__flag) begin
		if(ejection_channels_340__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_340__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_339__flag) begin
		if(ejection_channels_339__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_339__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_338__flag) begin
		if(ejection_channels_338__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_338__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_337__flag) begin
		if(ejection_channels_337__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_337__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_336__flag) begin
		if(ejection_channels_336__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_336__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_335__flag) begin
		if(ejection_channels_335__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_335__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_334__flag) begin
		if(ejection_channels_334__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_334__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_333__flag) begin
		if(ejection_channels_333__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_333__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_332__flag) begin
		if(ejection_channels_332__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_332__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_331__flag) begin
		if(ejection_channels_331__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_331__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_330__flag) begin
		if(ejection_channels_330__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_330__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_329__flag) begin
		if(ejection_channels_329__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_329__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_328__flag) begin
		if(ejection_channels_328__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_328__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_327__flag) begin
		if(ejection_channels_327__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_327__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_326__flag) begin
		if(ejection_channels_326__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_326__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_325__flag) begin
		if(ejection_channels_325__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_325__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_324__flag) begin
		if(ejection_channels_324__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_324__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_323__flag) begin
		if(ejection_channels_323__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_323__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_322__flag) begin
		if(ejection_channels_322__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_322__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_321__flag) begin
		if(ejection_channels_321__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_321__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_320__flag) begin
		if(ejection_channels_320__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_320__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_319__flag) begin
		if(ejection_channels_319__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_319__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_318__flag) begin
		if(ejection_channels_318__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_318__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_317__flag) begin
		if(ejection_channels_317__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_317__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_316__flag) begin
		if(ejection_channels_316__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_316__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_315__flag) begin
		if(ejection_channels_315__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_315__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_314__flag) begin
		if(ejection_channels_314__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_314__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_313__flag) begin
		if(ejection_channels_313__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_313__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_312__flag) begin
		if(ejection_channels_312__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_312__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_311__flag) begin
		if(ejection_channels_311__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_311__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_310__flag) begin
		if(ejection_channels_310__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_310__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_309__flag) begin
		if(ejection_channels_309__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_309__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_308__flag) begin
		if(ejection_channels_308__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_308__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_307__flag) begin
		if(ejection_channels_307__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_307__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_306__flag) begin
		if(ejection_channels_306__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_306__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_305__flag) begin
		if(ejection_channels_305__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_305__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_304__flag) begin
		if(ejection_channels_304__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_304__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_303__flag) begin
		if(ejection_channels_303__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_303__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_302__flag) begin
		if(ejection_channels_302__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_302__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_301__flag) begin
		if(ejection_channels_301__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_301__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_300__flag) begin
		if(ejection_channels_300__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_300__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_299__flag) begin
		if(ejection_channels_299__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_299__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_298__flag) begin
		if(ejection_channels_298__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_298__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_297__flag) begin
		if(ejection_channels_297__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_297__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_296__flag) begin
		if(ejection_channels_296__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_296__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_295__flag) begin
		if(ejection_channels_295__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_295__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_294__flag) begin
		if(ejection_channels_294__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_294__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_293__flag) begin
		if(ejection_channels_293__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_293__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_292__flag) begin
		if(ejection_channels_292__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_292__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_291__flag) begin
		if(ejection_channels_291__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_291__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_290__flag) begin
		if(ejection_channels_290__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_290__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_289__flag) begin
		if(ejection_channels_289__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_289__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_288__flag) begin
		if(ejection_channels_288__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_288__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_287__flag) begin
		if(ejection_channels_287__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_287__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_286__flag) begin
		if(ejection_channels_286__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_286__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_285__flag) begin
		if(ejection_channels_285__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_285__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_284__flag) begin
		if(ejection_channels_284__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_284__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_283__flag) begin
		if(ejection_channels_283__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_283__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_282__flag) begin
		if(ejection_channels_282__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_282__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_281__flag) begin
		if(ejection_channels_281__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_281__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_280__flag) begin
		if(ejection_channels_280__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_280__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_279__flag) begin
		if(ejection_channels_279__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_279__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_278__flag) begin
		if(ejection_channels_278__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_278__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_277__flag) begin
		if(ejection_channels_277__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_277__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_276__flag) begin
		if(ejection_channels_276__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_276__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_275__flag) begin
		if(ejection_channels_275__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_275__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_274__flag) begin
		if(ejection_channels_274__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_274__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_273__flag) begin
		if(ejection_channels_273__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_273__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_272__flag) begin
		if(ejection_channels_272__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_272__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_271__flag) begin
		if(ejection_channels_271__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_271__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_270__flag) begin
		if(ejection_channels_270__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_270__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_269__flag) begin
		if(ejection_channels_269__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_269__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_268__flag) begin
		if(ejection_channels_268__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_268__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_267__flag) begin
		if(ejection_channels_267__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_267__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_266__flag) begin
		if(ejection_channels_266__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_266__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_265__flag) begin
		if(ejection_channels_265__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_265__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_264__flag) begin
		if(ejection_channels_264__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_264__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_263__flag) begin
		if(ejection_channels_263__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_263__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_262__flag) begin
		if(ejection_channels_262__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_262__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_261__flag) begin
		if(ejection_channels_261__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_261__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_260__flag) begin
		if(ejection_channels_260__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_260__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_259__flag) begin
		if(ejection_channels_259__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_259__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_258__flag) begin
		if(ejection_channels_258__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_258__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_257__flag) begin
		if(ejection_channels_257__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_257__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_256__flag) begin
		if(ejection_channels_256__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_256__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_255__flag) begin
		if(ejection_channels_255__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_255__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_254__flag) begin
		if(ejection_channels_254__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_254__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_253__flag) begin
		if(ejection_channels_253__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_253__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_252__flag) begin
		if(ejection_channels_252__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_252__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_251__flag) begin
		if(ejection_channels_251__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_251__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_250__flag) begin
		if(ejection_channels_250__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_250__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_249__flag) begin
		if(ejection_channels_249__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_249__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_248__flag) begin
		if(ejection_channels_248__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_248__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_247__flag) begin
		if(ejection_channels_247__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_247__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_246__flag) begin
		if(ejection_channels_246__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_246__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_245__flag) begin
		if(ejection_channels_245__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_245__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_244__flag) begin
		if(ejection_channels_244__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_244__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_243__flag) begin
		if(ejection_channels_243__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_243__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_242__flag) begin
		if(ejection_channels_242__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_242__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_241__flag) begin
		if(ejection_channels_241__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_241__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_240__flag) begin
		if(ejection_channels_240__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_240__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_239__flag) begin
		if(ejection_channels_239__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_239__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_238__flag) begin
		if(ejection_channels_238__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_238__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_237__flag) begin
		if(ejection_channels_237__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_237__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_236__flag) begin
		if(ejection_channels_236__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_236__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_235__flag) begin
		if(ejection_channels_235__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_235__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_234__flag) begin
		if(ejection_channels_234__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_234__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_233__flag) begin
		if(ejection_channels_233__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_233__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_232__flag) begin
		if(ejection_channels_232__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_232__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_231__flag) begin
		if(ejection_channels_231__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_231__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_230__flag) begin
		if(ejection_channels_230__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_230__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_229__flag) begin
		if(ejection_channels_229__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_229__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_228__flag) begin
		if(ejection_channels_228__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_228__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_227__flag) begin
		if(ejection_channels_227__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_227__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_226__flag) begin
		if(ejection_channels_226__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_226__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_225__flag) begin
		if(ejection_channels_225__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_225__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_224__flag) begin
		if(ejection_channels_224__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_224__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_223__flag) begin
		if(ejection_channels_223__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_223__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_222__flag) begin
		if(ejection_channels_222__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_222__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_221__flag) begin
		if(ejection_channels_221__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_221__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_220__flag) begin
		if(ejection_channels_220__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_220__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_219__flag) begin
		if(ejection_channels_219__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_219__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_218__flag) begin
		if(ejection_channels_218__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_218__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_217__flag) begin
		if(ejection_channels_217__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_217__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_216__flag) begin
		if(ejection_channels_216__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_216__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_215__flag) begin
		if(ejection_channels_215__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_215__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_214__flag) begin
		if(ejection_channels_214__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_214__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_213__flag) begin
		if(ejection_channels_213__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_213__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_212__flag) begin
		if(ejection_channels_212__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_212__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_211__flag) begin
		if(ejection_channels_211__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_211__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_210__flag) begin
		if(ejection_channels_210__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_210__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_209__flag) begin
		if(ejection_channels_209__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_209__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_208__flag) begin
		if(ejection_channels_208__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_208__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_207__flag) begin
		if(ejection_channels_207__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_207__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_206__flag) begin
		if(ejection_channels_206__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_206__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_205__flag) begin
		if(ejection_channels_205__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_205__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_204__flag) begin
		if(ejection_channels_204__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_204__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_203__flag) begin
		if(ejection_channels_203__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_203__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_202__flag) begin
		if(ejection_channels_202__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_202__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_201__flag) begin
		if(ejection_channels_201__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_201__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_200__flag) begin
		if(ejection_channels_200__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_200__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_199__flag) begin
		if(ejection_channels_199__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_199__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_198__flag) begin
		if(ejection_channels_198__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_198__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_197__flag) begin
		if(ejection_channels_197__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_197__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_196__flag) begin
		if(ejection_channels_196__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_196__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_195__flag) begin
		if(ejection_channels_195__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_195__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_194__flag) begin
		if(ejection_channels_194__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_194__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_193__flag) begin
		if(ejection_channels_193__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_193__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_192__flag) begin
		if(ejection_channels_192__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_192__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_191__flag) begin
		if(ejection_channels_191__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_191__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_190__flag) begin
		if(ejection_channels_190__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_190__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_189__flag) begin
		if(ejection_channels_189__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_189__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_188__flag) begin
		if(ejection_channels_188__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_188__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_187__flag) begin
		if(ejection_channels_187__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_187__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_186__flag) begin
		if(ejection_channels_186__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_186__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_185__flag) begin
		if(ejection_channels_185__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_185__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_184__flag) begin
		if(ejection_channels_184__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_184__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_183__flag) begin
		if(ejection_channels_183__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_183__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_182__flag) begin
		if(ejection_channels_182__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_182__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_181__flag) begin
		if(ejection_channels_181__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_181__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_180__flag) begin
		if(ejection_channels_180__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_180__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_179__flag) begin
		if(ejection_channels_179__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_179__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_178__flag) begin
		if(ejection_channels_178__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_178__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_177__flag) begin
		if(ejection_channels_177__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_177__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_176__flag) begin
		if(ejection_channels_176__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_176__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_175__flag) begin
		if(ejection_channels_175__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_175__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_174__flag) begin
		if(ejection_channels_174__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_174__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_173__flag) begin
		if(ejection_channels_173__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_173__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_172__flag) begin
		if(ejection_channels_172__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_172__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_171__flag) begin
		if(ejection_channels_171__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_171__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_170__flag) begin
		if(ejection_channels_170__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_170__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_169__flag) begin
		if(ejection_channels_169__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_169__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_168__flag) begin
		if(ejection_channels_168__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_168__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_167__flag) begin
		if(ejection_channels_167__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_167__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_166__flag) begin
		if(ejection_channels_166__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_166__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_165__flag) begin
		if(ejection_channels_165__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_165__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_164__flag) begin
		if(ejection_channels_164__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_164__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_163__flag) begin
		if(ejection_channels_163__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_163__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_162__flag) begin
		if(ejection_channels_162__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_162__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_161__flag) begin
		if(ejection_channels_161__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_161__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_160__flag) begin
		if(ejection_channels_160__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_160__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_159__flag) begin
		if(ejection_channels_159__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_159__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_158__flag) begin
		if(ejection_channels_158__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_158__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_157__flag) begin
		if(ejection_channels_157__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_157__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_156__flag) begin
		if(ejection_channels_156__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_156__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_155__flag) begin
		if(ejection_channels_155__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_155__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_154__flag) begin
		if(ejection_channels_154__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_154__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_153__flag) begin
		if(ejection_channels_153__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_153__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_152__flag) begin
		if(ejection_channels_152__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_152__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_151__flag) begin
		if(ejection_channels_151__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_151__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_150__flag) begin
		if(ejection_channels_150__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_150__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_149__flag) begin
		if(ejection_channels_149__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_149__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_148__flag) begin
		if(ejection_channels_148__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_148__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_147__flag) begin
		if(ejection_channels_147__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_147__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_146__flag) begin
		if(ejection_channels_146__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_146__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_145__flag) begin
		if(ejection_channels_145__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_145__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_144__flag) begin
		if(ejection_channels_144__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_144__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_143__flag) begin
		if(ejection_channels_143__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_143__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_142__flag) begin
		if(ejection_channels_142__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_142__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_141__flag) begin
		if(ejection_channels_141__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_141__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_140__flag) begin
		if(ejection_channels_140__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_140__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_139__flag) begin
		if(ejection_channels_139__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_139__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_138__flag) begin
		if(ejection_channels_138__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_138__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_137__flag) begin
		if(ejection_channels_137__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_137__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_136__flag) begin
		if(ejection_channels_136__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_136__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_135__flag) begin
		if(ejection_channels_135__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_135__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_134__flag) begin
		if(ejection_channels_134__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_134__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_133__flag) begin
		if(ejection_channels_133__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_133__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_132__flag) begin
		if(ejection_channels_132__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_132__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_131__flag) begin
		if(ejection_channels_131__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_131__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_130__flag) begin
		if(ejection_channels_130__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_130__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_129__flag) begin
		if(ejection_channels_129__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_129__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_128__flag) begin
		if(ejection_channels_128__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_128__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_127__flag) begin
		if(ejection_channels_127__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_127__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_126__flag) begin
		if(ejection_channels_126__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_126__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_125__flag) begin
		if(ejection_channels_125__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_125__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_124__flag) begin
		if(ejection_channels_124__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_124__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_123__flag) begin
		if(ejection_channels_123__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_123__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_122__flag) begin
		if(ejection_channels_122__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_122__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_121__flag) begin
		if(ejection_channels_121__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_121__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_120__flag) begin
		if(ejection_channels_120__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_120__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_119__flag) begin
		if(ejection_channels_119__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_119__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_118__flag) begin
		if(ejection_channels_118__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_118__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_117__flag) begin
		if(ejection_channels_117__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_117__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_116__flag) begin
		if(ejection_channels_116__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_116__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_115__flag) begin
		if(ejection_channels_115__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_115__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_114__flag) begin
		if(ejection_channels_114__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_114__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_113__flag) begin
		if(ejection_channels_113__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_113__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_112__flag) begin
		if(ejection_channels_112__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_112__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_111__flag) begin
		if(ejection_channels_111__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_111__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_110__flag) begin
		if(ejection_channels_110__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_110__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_109__flag) begin
		if(ejection_channels_109__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_109__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_108__flag) begin
		if(ejection_channels_108__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_108__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_107__flag) begin
		if(ejection_channels_107__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_107__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_106__flag) begin
		if(ejection_channels_106__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_106__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_105__flag) begin
		if(ejection_channels_105__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_105__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_104__flag) begin
		if(ejection_channels_104__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_104__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_103__flag) begin
		if(ejection_channels_103__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_103__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_102__flag) begin
		if(ejection_channels_102__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_102__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_101__flag) begin
		if(ejection_channels_101__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_101__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_100__flag) begin
		if(ejection_channels_100__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_100__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_99__flag) begin
		if(ejection_channels_99__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_99__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_98__flag) begin
		if(ejection_channels_98__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_98__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_97__flag) begin
		if(ejection_channels_97__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_97__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_96__flag) begin
		if(ejection_channels_96__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_96__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_95__flag) begin
		if(ejection_channels_95__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_95__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_94__flag) begin
		if(ejection_channels_94__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_94__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_93__flag) begin
		if(ejection_channels_93__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_93__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_92__flag) begin
		if(ejection_channels_92__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_92__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_91__flag) begin
		if(ejection_channels_91__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_91__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_90__flag) begin
		if(ejection_channels_90__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_90__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_89__flag) begin
		if(ejection_channels_89__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_89__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_88__flag) begin
		if(ejection_channels_88__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_88__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_87__flag) begin
		if(ejection_channels_87__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_87__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_86__flag) begin
		if(ejection_channels_86__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_86__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_85__flag) begin
		if(ejection_channels_85__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_85__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_84__flag) begin
		if(ejection_channels_84__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_84__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_83__flag) begin
		if(ejection_channels_83__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_83__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_82__flag) begin
		if(ejection_channels_82__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_82__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_81__flag) begin
		if(ejection_channels_81__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_81__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_80__flag) begin
		if(ejection_channels_80__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_80__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_79__flag) begin
		if(ejection_channels_79__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_79__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_78__flag) begin
		if(ejection_channels_78__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_78__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_77__flag) begin
		if(ejection_channels_77__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_77__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_76__flag) begin
		if(ejection_channels_76__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_76__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_75__flag) begin
		if(ejection_channels_75__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_75__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_74__flag) begin
		if(ejection_channels_74__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_74__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_73__flag) begin
		if(ejection_channels_73__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_73__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_72__flag) begin
		if(ejection_channels_72__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_72__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_71__flag) begin
		if(ejection_channels_71__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_71__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_70__flag) begin
		if(ejection_channels_70__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_70__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_69__flag) begin
		if(ejection_channels_69__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_69__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_68__flag) begin
		if(ejection_channels_68__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_68__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_67__flag) begin
		if(ejection_channels_67__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_67__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_66__flag) begin
		if(ejection_channels_66__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_66__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_65__flag) begin
		if(ejection_channels_65__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_65__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_64__flag) begin
		if(ejection_channels_64__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_64__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_63__flag) begin
		if(ejection_channels_63__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_63__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_62__flag) begin
		if(ejection_channels_62__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_62__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_61__flag) begin
		if(ejection_channels_61__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_61__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_60__flag) begin
		if(ejection_channels_60__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_60__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_59__flag) begin
		if(ejection_channels_59__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_59__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_58__flag) begin
		if(ejection_channels_58__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_58__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_57__flag) begin
		if(ejection_channels_57__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_57__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_56__flag) begin
		if(ejection_channels_56__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_56__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_55__flag) begin
		if(ejection_channels_55__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_55__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_54__flag) begin
		if(ejection_channels_54__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_54__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_53__flag) begin
		if(ejection_channels_53__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_53__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_52__flag) begin
		if(ejection_channels_52__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_52__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_51__flag) begin
		if(ejection_channels_51__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_51__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_50__flag) begin
		if(ejection_channels_50__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_50__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_49__flag) begin
		if(ejection_channels_49__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_49__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_48__flag) begin
		if(ejection_channels_48__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_48__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_47__flag) begin
		if(ejection_channels_47__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_47__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_46__flag) begin
		if(ejection_channels_46__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_46__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_45__flag) begin
		if(ejection_channels_45__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_45__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_44__flag) begin
		if(ejection_channels_44__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_44__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_43__flag) begin
		if(ejection_channels_43__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_43__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_42__flag) begin
		if(ejection_channels_42__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_42__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_41__flag) begin
		if(ejection_channels_41__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_41__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_40__flag) begin
		if(ejection_channels_40__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_40__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_39__flag) begin
		if(ejection_channels_39__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_39__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_38__flag) begin
		if(ejection_channels_38__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_38__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_37__flag) begin
		if(ejection_channels_37__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_37__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_36__flag) begin
		if(ejection_channels_36__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_36__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_35__flag) begin
		if(ejection_channels_35__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_35__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_34__flag) begin
		if(ejection_channels_34__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_34__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_33__flag) begin
		if(ejection_channels_33__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_33__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_32__flag) begin
		if(ejection_channels_32__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_32__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_31__flag) begin
		if(ejection_channels_31__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_31__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_30__flag) begin
		if(ejection_channels_30__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_30__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_29__flag) begin
		if(ejection_channels_29__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_29__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_28__flag) begin
		if(ejection_channels_28__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_28__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_27__flag) begin
		if(ejection_channels_27__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_27__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_26__flag) begin
		if(ejection_channels_26__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_26__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_25__flag) begin
		if(ejection_channels_25__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_25__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_24__flag) begin
		if(ejection_channels_24__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_24__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_23__flag) begin
		if(ejection_channels_23__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_23__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_22__flag) begin
		if(ejection_channels_22__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_22__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_21__flag) begin
		if(ejection_channels_21__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_21__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_20__flag) begin
		if(ejection_channels_20__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_20__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_19__flag) begin
		if(ejection_channels_19__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_19__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_18__flag) begin
		if(ejection_channels_18__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_18__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_17__flag) begin
		if(ejection_channels_17__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_17__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_16__flag) begin
		if(ejection_channels_16__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_16__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_15__flag) begin
		if(ejection_channels_15__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_15__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_14__flag) begin
		if(ejection_channels_14__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_14__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_13__flag) begin
		if(ejection_channels_13__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_13__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_12__flag) begin
		if(ejection_channels_12__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_12__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_11__flag) begin
		if(ejection_channels_11__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_11__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_10__flag) begin
		if(ejection_channels_10__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_10__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_9__flag) begin
		if(ejection_channels_9__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_9__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_8__flag) begin
		if(ejection_channels_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_7__flag) begin
		if(ejection_channels_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_6__flag) begin
		if(ejection_channels_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_5__flag) begin
		if(ejection_channels_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_4__flag) begin
		if(ejection_channels_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_3__flag) begin
		if(ejection_channels_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_2__flag) begin
		if(ejection_channels_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_1__flag) begin
		if(ejection_channels_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge ejection_channels_0__flag) begin
		if(ejection_channels_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on ejection_channels_0__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_8__flag) begin
		if(rtr_error_8__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_8__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_7__flag) begin
		if(rtr_error_7__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_7__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_6__flag) begin
		if(rtr_error_6__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_6__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_5__flag) begin
		if(rtr_error_5__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_5__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_4__flag) begin
		if(rtr_error_4__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_4__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_3__flag) begin
		if(rtr_error_3__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_3__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_2__flag) begin
		if(rtr_error_2__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_2__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_1__flag) begin
		if(rtr_error_1__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_1__gfpga at time = %t", $realtime);
		end
	end

	always@(posedge rtr_error_0__flag) begin
		if(rtr_error_0__flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on rtr_error_0__gfpga at time = %t", $realtime);
		end
	end


// ----- Begin output waveform to VCD file-------
	initial begin
		$dumpfile("router_mesh_formal.vcd");
		$dumpvars(1, router_mesh_top_formal_verification_random_tb);
	end
// ----- END output waveform to VCD file -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#20
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for router_mesh_top_formal_verification_random_tb -----

