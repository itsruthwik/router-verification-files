//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[1][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Jun 27 10:27:38 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_1__2_ -----
module sb_1__2_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:188] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:188] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:188] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_;
//----- INPUT PORTS -----
input [0:188] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:188] chany_top_out;
//----- OUTPUT PORTS -----
output [0:188] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:188] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:188] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:4] mux_tree_tapbuf_size17_0_sram;
wire [0:4] mux_tree_tapbuf_size17_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size17_mem_0_ccff_tail;
wire [0:4] mux_tree_tapbuf_size18_0_sram;
wire [0:4] mux_tree_tapbuf_size18_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_10_sram;
wire [0:4] mux_tree_tapbuf_size18_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_11_sram;
wire [0:4] mux_tree_tapbuf_size18_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_12_sram;
wire [0:4] mux_tree_tapbuf_size18_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_13_sram;
wire [0:4] mux_tree_tapbuf_size18_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_14_sram;
wire [0:4] mux_tree_tapbuf_size18_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_15_sram;
wire [0:4] mux_tree_tapbuf_size18_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_1_sram;
wire [0:4] mux_tree_tapbuf_size18_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_2_sram;
wire [0:4] mux_tree_tapbuf_size18_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_3_sram;
wire [0:4] mux_tree_tapbuf_size18_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_4_sram;
wire [0:4] mux_tree_tapbuf_size18_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_5_sram;
wire [0:4] mux_tree_tapbuf_size18_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_6_sram;
wire [0:4] mux_tree_tapbuf_size18_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_7_sram;
wire [0:4] mux_tree_tapbuf_size18_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_8_sram;
wire [0:4] mux_tree_tapbuf_size18_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size18_9_sram;
wire [0:4] mux_tree_tapbuf_size18_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size18_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size18_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size19_0_sram;
wire [0:4] mux_tree_tapbuf_size19_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_10_sram;
wire [0:4] mux_tree_tapbuf_size19_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_11_sram;
wire [0:4] mux_tree_tapbuf_size19_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_12_sram;
wire [0:4] mux_tree_tapbuf_size19_12_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_13_sram;
wire [0:4] mux_tree_tapbuf_size19_13_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_14_sram;
wire [0:4] mux_tree_tapbuf_size19_14_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_15_sram;
wire [0:4] mux_tree_tapbuf_size19_15_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_16_sram;
wire [0:4] mux_tree_tapbuf_size19_16_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_17_sram;
wire [0:4] mux_tree_tapbuf_size19_17_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_18_sram;
wire [0:4] mux_tree_tapbuf_size19_18_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_19_sram;
wire [0:4] mux_tree_tapbuf_size19_19_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_1_sram;
wire [0:4] mux_tree_tapbuf_size19_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_20_sram;
wire [0:4] mux_tree_tapbuf_size19_20_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_21_sram;
wire [0:4] mux_tree_tapbuf_size19_21_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_22_sram;
wire [0:4] mux_tree_tapbuf_size19_22_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_23_sram;
wire [0:4] mux_tree_tapbuf_size19_23_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_24_sram;
wire [0:4] mux_tree_tapbuf_size19_24_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_25_sram;
wire [0:4] mux_tree_tapbuf_size19_25_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_26_sram;
wire [0:4] mux_tree_tapbuf_size19_26_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_27_sram;
wire [0:4] mux_tree_tapbuf_size19_27_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_28_sram;
wire [0:4] mux_tree_tapbuf_size19_28_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_29_sram;
wire [0:4] mux_tree_tapbuf_size19_29_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_2_sram;
wire [0:4] mux_tree_tapbuf_size19_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_30_sram;
wire [0:4] mux_tree_tapbuf_size19_30_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_31_sram;
wire [0:4] mux_tree_tapbuf_size19_31_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_32_sram;
wire [0:4] mux_tree_tapbuf_size19_32_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_33_sram;
wire [0:4] mux_tree_tapbuf_size19_33_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_34_sram;
wire [0:4] mux_tree_tapbuf_size19_34_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_35_sram;
wire [0:4] mux_tree_tapbuf_size19_35_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_36_sram;
wire [0:4] mux_tree_tapbuf_size19_36_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_37_sram;
wire [0:4] mux_tree_tapbuf_size19_37_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_38_sram;
wire [0:4] mux_tree_tapbuf_size19_38_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_39_sram;
wire [0:4] mux_tree_tapbuf_size19_39_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_3_sram;
wire [0:4] mux_tree_tapbuf_size19_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_40_sram;
wire [0:4] mux_tree_tapbuf_size19_40_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_41_sram;
wire [0:4] mux_tree_tapbuf_size19_41_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_42_sram;
wire [0:4] mux_tree_tapbuf_size19_42_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_43_sram;
wire [0:4] mux_tree_tapbuf_size19_43_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_44_sram;
wire [0:4] mux_tree_tapbuf_size19_44_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_45_sram;
wire [0:4] mux_tree_tapbuf_size19_45_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_46_sram;
wire [0:4] mux_tree_tapbuf_size19_46_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_47_sram;
wire [0:4] mux_tree_tapbuf_size19_47_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_48_sram;
wire [0:4] mux_tree_tapbuf_size19_48_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_49_sram;
wire [0:4] mux_tree_tapbuf_size19_49_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_4_sram;
wire [0:4] mux_tree_tapbuf_size19_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_50_sram;
wire [0:4] mux_tree_tapbuf_size19_50_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_51_sram;
wire [0:4] mux_tree_tapbuf_size19_51_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_52_sram;
wire [0:4] mux_tree_tapbuf_size19_52_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_53_sram;
wire [0:4] mux_tree_tapbuf_size19_53_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_54_sram;
wire [0:4] mux_tree_tapbuf_size19_54_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_55_sram;
wire [0:4] mux_tree_tapbuf_size19_55_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_56_sram;
wire [0:4] mux_tree_tapbuf_size19_56_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_57_sram;
wire [0:4] mux_tree_tapbuf_size19_57_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_58_sram;
wire [0:4] mux_tree_tapbuf_size19_58_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_59_sram;
wire [0:4] mux_tree_tapbuf_size19_59_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_5_sram;
wire [0:4] mux_tree_tapbuf_size19_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_60_sram;
wire [0:4] mux_tree_tapbuf_size19_60_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_61_sram;
wire [0:4] mux_tree_tapbuf_size19_61_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_62_sram;
wire [0:4] mux_tree_tapbuf_size19_62_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_63_sram;
wire [0:4] mux_tree_tapbuf_size19_63_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_64_sram;
wire [0:4] mux_tree_tapbuf_size19_64_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_65_sram;
wire [0:4] mux_tree_tapbuf_size19_65_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_66_sram;
wire [0:4] mux_tree_tapbuf_size19_66_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_6_sram;
wire [0:4] mux_tree_tapbuf_size19_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_7_sram;
wire [0:4] mux_tree_tapbuf_size19_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_8_sram;
wire [0:4] mux_tree_tapbuf_size19_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size19_9_sram;
wire [0:4] mux_tree_tapbuf_size19_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size19_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size19_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size20_0_sram;
wire [0:4] mux_tree_tapbuf_size20_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_10_sram;
wire [0:4] mux_tree_tapbuf_size20_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_11_sram;
wire [0:4] mux_tree_tapbuf_size20_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_1_sram;
wire [0:4] mux_tree_tapbuf_size20_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_2_sram;
wire [0:4] mux_tree_tapbuf_size20_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_3_sram;
wire [0:4] mux_tree_tapbuf_size20_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_4_sram;
wire [0:4] mux_tree_tapbuf_size20_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_5_sram;
wire [0:4] mux_tree_tapbuf_size20_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_6_sram;
wire [0:4] mux_tree_tapbuf_size20_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_7_sram;
wire [0:4] mux_tree_tapbuf_size20_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_8_sram;
wire [0:4] mux_tree_tapbuf_size20_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_9_sram;
wire [0:4] mux_tree_tapbuf_size20_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size20_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:3] mux_tree_tapbuf_size8_0_sram;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_10_sram;
wire [0:3] mux_tree_tapbuf_size8_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_11_sram;
wire [0:3] mux_tree_tapbuf_size8_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_12_sram;
wire [0:3] mux_tree_tapbuf_size8_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_13_sram;
wire [0:3] mux_tree_tapbuf_size8_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_14_sram;
wire [0:3] mux_tree_tapbuf_size8_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_15_sram;
wire [0:3] mux_tree_tapbuf_size8_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_16_sram;
wire [0:3] mux_tree_tapbuf_size8_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_17_sram;
wire [0:3] mux_tree_tapbuf_size8_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_18_sram;
wire [0:3] mux_tree_tapbuf_size8_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_19_sram;
wire [0:3] mux_tree_tapbuf_size8_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_1_sram;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_20_sram;
wire [0:3] mux_tree_tapbuf_size8_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_21_sram;
wire [0:3] mux_tree_tapbuf_size8_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_22_sram;
wire [0:3] mux_tree_tapbuf_size8_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_23_sram;
wire [0:3] mux_tree_tapbuf_size8_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_24_sram;
wire [0:3] mux_tree_tapbuf_size8_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_25_sram;
wire [0:3] mux_tree_tapbuf_size8_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_26_sram;
wire [0:3] mux_tree_tapbuf_size8_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_27_sram;
wire [0:3] mux_tree_tapbuf_size8_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_28_sram;
wire [0:3] mux_tree_tapbuf_size8_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_29_sram;
wire [0:3] mux_tree_tapbuf_size8_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_2_sram;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_30_sram;
wire [0:3] mux_tree_tapbuf_size8_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_31_sram;
wire [0:3] mux_tree_tapbuf_size8_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_32_sram;
wire [0:3] mux_tree_tapbuf_size8_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_33_sram;
wire [0:3] mux_tree_tapbuf_size8_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_34_sram;
wire [0:3] mux_tree_tapbuf_size8_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_35_sram;
wire [0:3] mux_tree_tapbuf_size8_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_36_sram;
wire [0:3] mux_tree_tapbuf_size8_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_37_sram;
wire [0:3] mux_tree_tapbuf_size8_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_38_sram;
wire [0:3] mux_tree_tapbuf_size8_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_39_sram;
wire [0:3] mux_tree_tapbuf_size8_39_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_3_sram;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_40_sram;
wire [0:3] mux_tree_tapbuf_size8_40_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_41_sram;
wire [0:3] mux_tree_tapbuf_size8_41_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_42_sram;
wire [0:3] mux_tree_tapbuf_size8_42_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_43_sram;
wire [0:3] mux_tree_tapbuf_size8_43_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_44_sram;
wire [0:3] mux_tree_tapbuf_size8_44_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_45_sram;
wire [0:3] mux_tree_tapbuf_size8_45_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_46_sram;
wire [0:3] mux_tree_tapbuf_size8_46_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_47_sram;
wire [0:3] mux_tree_tapbuf_size8_47_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_48_sram;
wire [0:3] mux_tree_tapbuf_size8_48_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_49_sram;
wire [0:3] mux_tree_tapbuf_size8_49_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_4_sram;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_50_sram;
wire [0:3] mux_tree_tapbuf_size8_50_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_51_sram;
wire [0:3] mux_tree_tapbuf_size8_51_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_52_sram;
wire [0:3] mux_tree_tapbuf_size8_52_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_53_sram;
wire [0:3] mux_tree_tapbuf_size8_53_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_54_sram;
wire [0:3] mux_tree_tapbuf_size8_54_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_55_sram;
wire [0:3] mux_tree_tapbuf_size8_55_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_56_sram;
wire [0:3] mux_tree_tapbuf_size8_56_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_57_sram;
wire [0:3] mux_tree_tapbuf_size8_57_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_58_sram;
wire [0:3] mux_tree_tapbuf_size8_58_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_59_sram;
wire [0:3] mux_tree_tapbuf_size8_59_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_5_sram;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_60_sram;
wire [0:3] mux_tree_tapbuf_size8_60_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_61_sram;
wire [0:3] mux_tree_tapbuf_size8_61_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_62_sram;
wire [0:3] mux_tree_tapbuf_size8_62_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_63_sram;
wire [0:3] mux_tree_tapbuf_size8_63_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_64_sram;
wire [0:3] mux_tree_tapbuf_size8_64_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_65_sram;
wire [0:3] mux_tree_tapbuf_size8_65_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_66_sram;
wire [0:3] mux_tree_tapbuf_size8_66_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_67_sram;
wire [0:3] mux_tree_tapbuf_size8_67_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_68_sram;
wire [0:3] mux_tree_tapbuf_size8_68_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_69_sram;
wire [0:3] mux_tree_tapbuf_size8_69_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_6_sram;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_70_sram;
wire [0:3] mux_tree_tapbuf_size8_70_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_71_sram;
wire [0:3] mux_tree_tapbuf_size8_71_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_72_sram;
wire [0:3] mux_tree_tapbuf_size8_72_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_7_sram;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_8_sram;
wire [0:3] mux_tree_tapbuf_size8_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_9_sram;
wire [0:3] mux_tree_tapbuf_size8_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_10_sram;
wire [0:3] mux_tree_tapbuf_size9_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_11_sram;
wire [0:3] mux_tree_tapbuf_size9_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_12_sram;
wire [0:3] mux_tree_tapbuf_size9_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_13_sram;
wire [0:3] mux_tree_tapbuf_size9_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_14_sram;
wire [0:3] mux_tree_tapbuf_size9_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_15_sram;
wire [0:3] mux_tree_tapbuf_size9_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_16_sram;
wire [0:3] mux_tree_tapbuf_size9_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_17_sram;
wire [0:3] mux_tree_tapbuf_size9_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_1_sram;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_2_sram;
wire [0:3] mux_tree_tapbuf_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_3_sram;
wire [0:3] mux_tree_tapbuf_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_4_sram;
wire [0:3] mux_tree_tapbuf_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_5_sram;
wire [0:3] mux_tree_tapbuf_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_6_sram;
wire [0:3] mux_tree_tapbuf_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_7_sram;
wire [0:3] mux_tree_tapbuf_size9_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_8_sram;
wire [0:3] mux_tree_tapbuf_size9_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_9_sram;
wire [0:3] mux_tree_tapbuf_size9_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[161] = chany_top_in[160];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[162] = chany_top_in[161];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[163] = chany_top_in[162];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[165] = chany_top_in[164];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[166] = chany_top_in[165];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[167] = chany_top_in[166];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[169] = chany_top_in[168];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[170] = chany_top_in[169];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[171] = chany_top_in[170];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[173] = chany_top_in[172];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[174] = chany_top_in[173];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[175] = chany_top_in[174];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[177] = chany_top_in[176];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[178] = chany_top_in[177];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[179] = chany_top_in[178];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[181] = chany_top_in[180];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[182] = chany_top_in[181];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[183] = chany_top_in[182];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[185] = chany_top_in[184];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[186] = chany_top_in[185];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[187] = chany_top_in[186];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[105] = chanx_right_in[104];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[106] = chanx_right_in[105];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[107] = chanx_right_in[106];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[109] = chanx_right_in[108];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[110] = chanx_right_in[109];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[111] = chanx_right_in[110];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[113] = chanx_right_in[112];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[114] = chanx_right_in[113];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[115] = chanx_right_in[114];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[117] = chanx_right_in[116];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[118] = chanx_right_in[117];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[119] = chanx_right_in[118];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[121] = chanx_right_in[120];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[122] = chanx_right_in[121];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[123] = chanx_right_in[122];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[125] = chanx_right_in[124];
// ----- Local connection due to Wire 316 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[126] = chanx_right_in[125];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[127] = chanx_right_in[126];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[129] = chanx_right_in[128];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[130] = chanx_right_in[129];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[131] = chanx_right_in[130];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[133] = chanx_right_in[132];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[134] = chanx_right_in[133];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[135] = chanx_right_in[134];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[137] = chanx_right_in[136];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[138] = chanx_right_in[137];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[139] = chanx_right_in[138];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[141] = chanx_right_in[140];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[142] = chanx_right_in[141];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[143] = chanx_right_in[142];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[145] = chanx_right_in[144];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[146] = chanx_right_in[145];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[147] = chanx_right_in[146];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[149] = chanx_right_in[148];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[150] = chanx_right_in[149];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[151] = chanx_right_in[150];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[153] = chanx_right_in[152];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[154] = chanx_right_in[153];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[155] = chanx_right_in[154];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[157] = chanx_right_in[156];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[158] = chanx_right_in[157];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[159] = chanx_right_in[158];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[161] = chanx_right_in[160];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[162] = chanx_right_in[161];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[163] = chanx_right_in[162];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[165] = chanx_right_in[164];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[166] = chanx_right_in[165];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[167] = chanx_right_in[166];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[169] = chanx_right_in[168];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[170] = chanx_right_in[169];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[171] = chanx_right_in[170];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[173] = chanx_right_in[172];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[174] = chanx_right_in[173];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[175] = chanx_right_in[174];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[177] = chanx_right_in[176];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[178] = chanx_right_in[177];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[179] = chanx_right_in[178];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[181] = chanx_right_in[180];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[182] = chanx_right_in[181];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[183] = chanx_right_in[182];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[185] = chanx_right_in[184];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[186] = chanx_right_in[185];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[187] = chanx_right_in[186];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 403 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 407 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 411 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 415 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 419 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 423 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 424 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 426 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 430 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 434 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 438 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 442 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 446 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 450 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 454 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 458 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 462 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 466 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 470 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 474 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 478 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 482 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 486 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 490 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 494 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 498 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 502 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 506 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 510 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 514 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 518 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 522 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 526 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 530 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 531 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 532 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 534 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 535 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 536 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 538 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 539 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 540 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- Local connection due to Wire 542 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[161] = chany_bottom_in[160];
// ----- Local connection due to Wire 543 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[162] = chany_bottom_in[161];
// ----- Local connection due to Wire 544 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[163] = chany_bottom_in[162];
// ----- Local connection due to Wire 546 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[165] = chany_bottom_in[164];
// ----- Local connection due to Wire 547 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[166] = chany_bottom_in[165];
// ----- Local connection due to Wire 548 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[167] = chany_bottom_in[166];
// ----- Local connection due to Wire 550 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[169] = chany_bottom_in[168];
// ----- Local connection due to Wire 551 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[170] = chany_bottom_in[169];
// ----- Local connection due to Wire 552 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[171] = chany_bottom_in[170];
// ----- Local connection due to Wire 554 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[173] = chany_bottom_in[172];
// ----- Local connection due to Wire 555 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[174] = chany_bottom_in[173];
// ----- Local connection due to Wire 556 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[175] = chany_bottom_in[174];
// ----- Local connection due to Wire 558 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[177] = chany_bottom_in[176];
// ----- Local connection due to Wire 559 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[178] = chany_bottom_in[177];
// ----- Local connection due to Wire 560 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[179] = chany_bottom_in[178];
// ----- Local connection due to Wire 562 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[181] = chany_bottom_in[180];
// ----- Local connection due to Wire 563 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[182] = chany_bottom_in[181];
// ----- Local connection due to Wire 564 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[183] = chany_bottom_in[182];
// ----- Local connection due to Wire 566 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[185] = chany_bottom_in[184];
// ----- Local connection due to Wire 567 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[186] = chany_bottom_in[185];
// ----- Local connection due to Wire 568 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[187] = chany_bottom_in[186];
// ----- Local connection due to Wire 660 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 661 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 662 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 664 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 665 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 666 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 668 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 669 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 670 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 672 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 673 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 674 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 676 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 677 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 678 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 680 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 681 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 682 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 684 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 685 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 686 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 688 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 689 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 690 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 692 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 693 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 694 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 696 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 697 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 698 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 700 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 701 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 702 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 704 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 705 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 706 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 708 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 709 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 710 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 712 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 713 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 714 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 716 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 717 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 718 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 720 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 721 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 722 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 724 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 725 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 726 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 728 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 729 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 730 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 732 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 733 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 734 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 736 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 737 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 738 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 740 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 741 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 742 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 744 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 745 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 746 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 748 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 749 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 750 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 752 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 753 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 754 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 756 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 757 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 758 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 760 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 761 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 762 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- Local connection due to Wire 764 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[105] = chanx_left_in[104];
// ----- Local connection due to Wire 765 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[106] = chanx_left_in[105];
// ----- Local connection due to Wire 766 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[107] = chanx_left_in[106];
// ----- Local connection due to Wire 768 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[109] = chanx_left_in[108];
// ----- Local connection due to Wire 769 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[110] = chanx_left_in[109];
// ----- Local connection due to Wire 770 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[111] = chanx_left_in[110];
// ----- Local connection due to Wire 772 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[113] = chanx_left_in[112];
// ----- Local connection due to Wire 773 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[114] = chanx_left_in[113];
// ----- Local connection due to Wire 774 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[115] = chanx_left_in[114];
// ----- Local connection due to Wire 776 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[117] = chanx_left_in[116];
// ----- Local connection due to Wire 777 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[118] = chanx_left_in[117];
// ----- Local connection due to Wire 778 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[119] = chanx_left_in[118];
// ----- Local connection due to Wire 780 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[121] = chanx_left_in[120];
// ----- Local connection due to Wire 781 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[122] = chanx_left_in[121];
// ----- Local connection due to Wire 782 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[123] = chanx_left_in[122];
// ----- Local connection due to Wire 784 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[125] = chanx_left_in[124];
// ----- Local connection due to Wire 785 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[126] = chanx_left_in[125];
// ----- Local connection due to Wire 786 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[127] = chanx_left_in[126];
// ----- Local connection due to Wire 788 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[129] = chanx_left_in[128];
// ----- Local connection due to Wire 789 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[130] = chanx_left_in[129];
// ----- Local connection due to Wire 790 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[131] = chanx_left_in[130];
// ----- Local connection due to Wire 792 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[133] = chanx_left_in[132];
// ----- Local connection due to Wire 793 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[134] = chanx_left_in[133];
// ----- Local connection due to Wire 794 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[135] = chanx_left_in[134];
// ----- Local connection due to Wire 796 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[137] = chanx_left_in[136];
// ----- Local connection due to Wire 797 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[138] = chanx_left_in[137];
// ----- Local connection due to Wire 798 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[139] = chanx_left_in[138];
// ----- Local connection due to Wire 800 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[141] = chanx_left_in[140];
// ----- Local connection due to Wire 801 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[142] = chanx_left_in[141];
// ----- Local connection due to Wire 802 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[143] = chanx_left_in[142];
// ----- Local connection due to Wire 804 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[145] = chanx_left_in[144];
// ----- Local connection due to Wire 805 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[146] = chanx_left_in[145];
// ----- Local connection due to Wire 806 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[147] = chanx_left_in[146];
// ----- Local connection due to Wire 808 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[149] = chanx_left_in[148];
// ----- Local connection due to Wire 809 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[150] = chanx_left_in[149];
// ----- Local connection due to Wire 810 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[151] = chanx_left_in[150];
// ----- Local connection due to Wire 812 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[153] = chanx_left_in[152];
// ----- Local connection due to Wire 813 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[154] = chanx_left_in[153];
// ----- Local connection due to Wire 814 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[155] = chanx_left_in[154];
// ----- Local connection due to Wire 816 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[157] = chanx_left_in[156];
// ----- Local connection due to Wire 817 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[158] = chanx_left_in[157];
// ----- Local connection due to Wire 818 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[159] = chanx_left_in[158];
// ----- Local connection due to Wire 820 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[161] = chanx_left_in[160];
// ----- Local connection due to Wire 821 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[162] = chanx_left_in[161];
// ----- Local connection due to Wire 822 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[163] = chanx_left_in[162];
// ----- Local connection due to Wire 824 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[165] = chanx_left_in[164];
// ----- Local connection due to Wire 825 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[166] = chanx_left_in[165];
// ----- Local connection due to Wire 826 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[167] = chanx_left_in[166];
// ----- Local connection due to Wire 828 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[169] = chanx_left_in[168];
// ----- Local connection due to Wire 829 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[170] = chanx_left_in[169];
// ----- Local connection due to Wire 830 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[171] = chanx_left_in[170];
// ----- Local connection due to Wire 832 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[173] = chanx_left_in[172];
// ----- Local connection due to Wire 833 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[174] = chanx_left_in[173];
// ----- Local connection due to Wire 834 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[175] = chanx_left_in[174];
// ----- Local connection due to Wire 836 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[177] = chanx_left_in[176];
// ----- Local connection due to Wire 837 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[178] = chanx_left_in[177];
// ----- Local connection due to Wire 838 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[179] = chanx_left_in[178];
// ----- Local connection due to Wire 840 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[181] = chanx_left_in[180];
// ----- Local connection due to Wire 841 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[182] = chanx_left_in[181];
// ----- Local connection due to Wire 842 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[183] = chanx_left_in[182];
// ----- Local connection due to Wire 844 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[185] = chanx_left_in[184];
// ----- Local connection due to Wire 845 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[186] = chanx_left_in[185];
// ----- Local connection due to Wire 846 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[187] = chanx_left_in[186];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size9 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[65], chanx_right_in[129], chanx_left_in[0], chanx_left_in[3], chanx_left_in[64], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size9 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[13], chanx_right_in[43], chanx_right_in[77], chanx_right_in[141], chanx_left_in[52], chanx_left_in[116], chanx_left_in[159], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_1_sram_inv[0:3]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size9 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[14], chanx_right_in[47], chanx_right_in[78], chanx_right_in[142], chanx_left_in[50], chanx_left_in[114], chanx_left_in[155], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_2_sram_inv[0:3]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size9 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[25], chanx_right_in[79], chanx_right_in[89], chanx_right_in[153], chanx_left_in[40], chanx_left_in[104], chanx_left_in[123], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_3_sram_inv[0:3]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size9 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[26], chanx_right_in[83], chanx_right_in[90], chanx_right_in[154], chanx_left_in[38], chanx_left_in[102], chanx_left_in[119], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_4_sram_inv[0:3]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size9 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[37], chanx_right_in[101], chanx_right_in[115], chanx_right_in[165], chanx_left_in[28], chanx_left_in[87], chanx_left_in[92], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_5_sram_inv[0:3]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size9 mux_top_track_224 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[38], chanx_right_in[102], chanx_right_in[119], chanx_right_in[166], chanx_left_in[26], chanx_left_in[83], chanx_left_in[90], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_6_sram_inv[0:3]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size9 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[49], chanx_right_in[113], chanx_right_in[151], chanx_right_in[177], chanx_left_in[16], chanx_left_in[51], chanx_left_in[80], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_7_sram_inv[0:3]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size9 mux_top_track_296 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[50], chanx_right_in[114], chanx_right_in[155], chanx_right_in[178], chanx_left_in[14], chanx_left_in[47], chanx_left_in[78], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size9_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_8_sram_inv[0:3]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size9 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[74], chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[49], chany_bottom_in[113], chany_bottom_in[151], chany_bottom_in[177]}),
		.sram(mux_tree_tapbuf_size9_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_9_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size9 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[76], chany_top_in[140], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[48], chany_bottom_in[112], chany_bottom_in[147], chany_bottom_in[176]}),
		.sram(mux_tree_tapbuf_size9_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_10_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size9 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[86], chany_top_in[150], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[37], chany_bottom_in[101], chany_bottom_in[115], chany_bottom_in[165]}),
		.sram(mux_tree_tapbuf_size9_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_11_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size9 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[88], chany_top_in[152], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[36], chany_bottom_in[100], chany_bottom_in[111], chany_bottom_in[164]}),
		.sram(mux_tree_tapbuf_size9_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_12_sram_inv[0:3]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size9 mux_right_track_216 (
		.in({chany_top_in[34], chany_top_in[98], chany_top_in[107], chany_top_in[162], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[89], chany_bottom_in[153]}),
		.sram(mux_tree_tapbuf_size9_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_13_sram_inv[0:3]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size9 mux_right_track_224 (
		.in({chany_top_in[36], chany_top_in[100], chany_top_in[111], chany_top_in[164], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[88], chany_bottom_in[152]}),
		.sram(mux_tree_tapbuf_size9_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_14_sram_inv[0:3]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size9 mux_right_track_288 (
		.in({chany_top_in[46], chany_top_in[110], chany_top_in[143], chany_top_in[174], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[77], chany_bottom_in[141]}),
		.sram(mux_tree_tapbuf_size9_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_15_sram_inv[0:3]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size9 mux_right_track_296 (
		.in({chany_top_in[48], chany_top_in[112], chany_top_in[147], chany_top_in[176], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[76], chany_bottom_in[140]}),
		.sram(mux_tree_tapbuf_size9_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_16_sram_inv[0:3]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size9 mux_right_track_360 (
		.in({chany_top_in[58], chany_top_in[122], chany_top_in[179], chany_top_in[186], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[65], chany_bottom_in[129]}),
		.sram(mux_tree_tapbuf_size9_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_17_sram_inv[0:3]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size9_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_8_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_9_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_10_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_11_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_12_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_13_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_14_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_15_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_16_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_17_sram_inv[0:3]));

	mux_tree_tapbuf_size8 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[66], chanx_right_in[130], chanx_left_in[62], chanx_left_in[126], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size8_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_0_sram_inv[0:3]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size8 mux_top_track_32 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[70], chanx_right_in[134], chanx_left_in[58], chanx_left_in[122], chanx_left_in[179], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size8_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_1_sram_inv[0:3]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size8 mux_top_track_40 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[72], chanx_right_in[136], chanx_left_in[57], chanx_left_in[121], chanx_left_in[175], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size8_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_2_sram_inv[0:3]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size8 mux_top_track_48 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[73], chanx_right_in[137], chanx_left_in[56], chanx_left_in[120], chanx_left_in[171], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size8_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_3_sram_inv[0:3]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size8 mux_top_track_56 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[74], chanx_right_in[138], chanx_left_in[54], chanx_left_in[118], chanx_left_in[167], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size8_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_4_sram_inv[0:3]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size8 mux_top_track_64 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[76], chanx_right_in[140], chanx_left_in[53], chanx_left_in[117], chanx_left_in[163], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size8_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_5_sram_inv[0:3]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size8 mux_top_track_88 (
		.in({chanx_right_in[16], chanx_right_in[51], chanx_right_in[80], chanx_right_in[144], chanx_left_in[49], chanx_left_in[113], chanx_left_in[151], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size8_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_6_sram_inv[0:3]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size8 mux_top_track_96 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[81], chanx_right_in[145], chanx_left_in[48], chanx_left_in[112], chanx_left_in[147], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size8_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_7_sram_inv[0:3]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size8 mux_top_track_104 (
		.in({chanx_right_in[18], chanx_right_in[59], chanx_right_in[82], chanx_right_in[146], chanx_left_in[46], chanx_left_in[110], chanx_left_in[143], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size8_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_8_sram_inv[0:3]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size8 mux_top_track_112 (
		.in({chanx_right_in[20], chanx_right_in[63], chanx_right_in[84], chanx_right_in[148], chanx_left_in[45], chanx_left_in[109], chanx_left_in[139], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size8_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_9_sram_inv[0:3]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size8 mux_top_track_120 (
		.in({chanx_right_in[21], chanx_right_in[67], chanx_right_in[85], chanx_right_in[149], chanx_left_in[44], chanx_left_in[108], chanx_left_in[135], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size8_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_10_sram_inv[0:3]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size8 mux_top_track_128 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[86], chanx_right_in[150], chanx_left_in[42], chanx_left_in[106], chanx_left_in[131], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size8_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_11_sram_inv[0:3]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size8 mux_top_track_136 (
		.in({chanx_right_in[24], chanx_right_in[75], chanx_right_in[88], chanx_right_in[152], chanx_left_in[41], chanx_left_in[105], chanx_left_in[127], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size8_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_12_sram_inv[0:3]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size8 mux_top_track_160 (
		.in({chanx_right_in[28], chanx_right_in[87], chanx_right_in[92], chanx_right_in[156], chanx_left_in[37], chanx_left_in[101], chanx_left_in[115], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size8_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_13_sram_inv[0:3]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size8 mux_top_track_168 (
		.in({chanx_right_in[29], chanx_right_in[91], chanx_right_in[93], chanx_right_in[157], chanx_left_in[36], chanx_left_in[100], chanx_left_in[111], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size8_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_14_sram_inv[0:3]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size8 mux_top_track_176 (
		.in({chanx_right_in[30], chanx_right_in[94:95], chanx_right_in[158], chanx_left_in[34], chanx_left_in[98], chanx_left_in[107], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size8_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_15_sram_inv[0:3]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size8 mux_top_track_184 (
		.in({chanx_right_in[32], chanx_right_in[96], chanx_right_in[99], chanx_right_in[160], chanx_left_in[33], chanx_left_in[97], chanx_left_in[103], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size8_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_16_sram_inv[0:3]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size8 mux_top_track_192 (
		.in({chanx_right_in[33], chanx_right_in[97], chanx_right_in[103], chanx_right_in[161], chanx_left_in[32], chanx_left_in[96], chanx_left_in[99], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size8_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_17_sram_inv[0:3]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size8 mux_top_track_200 (
		.in({chanx_right_in[34], chanx_right_in[98], chanx_right_in[107], chanx_right_in[162], chanx_left_in[30], chanx_left_in[94:95], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size8_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_18_sram_inv[0:3]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size8 mux_top_track_208 (
		.in({chanx_right_in[36], chanx_right_in[100], chanx_right_in[111], chanx_right_in[164], chanx_left_in[29], chanx_left_in[91], chanx_left_in[93], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size8_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_19_sram_inv[0:3]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size8 mux_top_track_232 (
		.in({chanx_right_in[40], chanx_right_in[104], chanx_right_in[123], chanx_right_in[168], chanx_left_in[25], chanx_left_in[79], chanx_left_in[89], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size8_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_20_sram_inv[0:3]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size8 mux_top_track_240 (
		.in({chanx_right_in[41], chanx_right_in[105], chanx_right_in[127], chanx_right_in[169], chanx_left_in[24], chanx_left_in[75], chanx_left_in[88], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size8_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_21_sram_inv[0:3]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size8 mux_top_track_248 (
		.in({chanx_right_in[42], chanx_right_in[106], chanx_right_in[131], chanx_right_in[170], chanx_left_in[22], chanx_left_in[71], chanx_left_in[86], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size8_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_22_sram_inv[0:3]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size8 mux_top_track_256 (
		.in({chanx_right_in[44], chanx_right_in[108], chanx_right_in[135], chanx_right_in[172], chanx_left_in[21], chanx_left_in[67], chanx_left_in[85], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size8_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_23_sram_inv[0:3]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size8 mux_top_track_264 (
		.in({chanx_right_in[45], chanx_right_in[109], chanx_right_in[139], chanx_right_in[173], chanx_left_in[20], chanx_left_in[63], chanx_left_in[84], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size8_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_24_sram_inv[0:3]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size8 mux_top_track_272 (
		.in({chanx_right_in[46], chanx_right_in[110], chanx_right_in[143], chanx_right_in[174], chanx_left_in[18], chanx_left_in[59], chanx_left_in[82], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size8_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_25_sram_inv[0:3]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size8 mux_top_track_280 (
		.in({chanx_right_in[48], chanx_right_in[112], chanx_right_in[147], chanx_right_in[176], chanx_left_in[17], chanx_left_in[55], chanx_left_in[81], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size8_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_26_sram_inv[0:3]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size8 mux_top_track_304 (
		.in({chanx_right_in[52], chanx_right_in[116], chanx_right_in[159], chanx_right_in[180], chanx_left_in[13], chanx_left_in[43], chanx_left_in[77], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size8_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_27_sram_inv[0:3]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size8 mux_top_track_312 (
		.in({chanx_right_in[53], chanx_right_in[117], chanx_right_in[163], chanx_right_in[181], chanx_left_in[12], chanx_left_in[39], chanx_left_in[76], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size8_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_28_sram_inv[0:3]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size8 mux_top_track_320 (
		.in({chanx_right_in[54], chanx_right_in[118], chanx_right_in[167], chanx_right_in[182], chanx_left_in[10], chanx_left_in[35], chanx_left_in[74], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size8_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_29_sram_inv[0:3]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size8 mux_top_track_328 (
		.in({chanx_right_in[56], chanx_right_in[120], chanx_right_in[171], chanx_right_in[184], chanx_left_in[9], chanx_left_in[31], chanx_left_in[73], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size8_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_30_sram_inv[0:3]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size8 mux_top_track_336 (
		.in({chanx_right_in[57], chanx_right_in[121], chanx_right_in[175], chanx_right_in[185], chanx_left_in[8], chanx_left_in[27], chanx_left_in[72], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size8_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_31_sram_inv[0:3]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size8 mux_top_track_344 (
		.in({chanx_right_in[58], chanx_right_in[122], chanx_right_in[179], chanx_right_in[186], chanx_left_in[6], chanx_left_in[23], chanx_left_in[70], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size8_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_32_sram_inv[0:3]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size8 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_right_in[61], chanx_right_in[125], chanx_right_in[187], chanx_left_in[4], chanx_left_in[15], chanx_left_in[68], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size8_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_33_sram_inv[0:3]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size8 mux_top_track_368 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[62], chanx_right_in[126], chanx_right_in[188], chanx_left_in[2], chanx_left_in[11], chanx_left_in[66], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size8_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_34_sram_inv[0:3]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size8 mux_top_track_376 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[64], chanx_right_in[128], chanx_left_in[1], chanx_left_in[7], chanx_left_in[65], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size8_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_35_sram_inv[0:3]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size8 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[64], chany_top_in[128], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[60], chany_bottom_in[124], chany_bottom_in[183]}),
		.sram(mux_tree_tapbuf_size8_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_36_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size8 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[65], chany_top_in[129], chany_bottom_in[58], chany_bottom_in[122], chany_bottom_in[179], chany_bottom_in[186]}),
		.sram(mux_tree_tapbuf_size8_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_37_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size8 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[66], chany_top_in[130], chany_bottom_in[57], chany_bottom_in[121], chany_bottom_in[175], chany_bottom_in[185]}),
		.sram(mux_tree_tapbuf_size8_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_38_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size8 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[68], chany_top_in[132], chany_bottom_in[56], chany_bottom_in[120], chany_bottom_in[171], chany_bottom_in[184]}),
		.sram(mux_tree_tapbuf_size8_39_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_39_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size8 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[69], chany_top_in[133], chany_bottom_in[54], chany_bottom_in[118], chany_bottom_in[167], chany_bottom_in[182]}),
		.sram(mux_tree_tapbuf_size8_40_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_40_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size8 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[70], chany_top_in[134], chany_bottom_in[53], chany_bottom_in[117], chany_bottom_in[163], chany_bottom_in[181]}),
		.sram(mux_tree_tapbuf_size8_41_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_41_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size8 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[72], chany_top_in[136], chany_bottom_in[52], chany_bottom_in[116], chany_bottom_in[159], chany_bottom_in[180]}),
		.sram(mux_tree_tapbuf_size8_42_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_42_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size8 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[73], chany_top_in[137], chany_bottom_in[50], chany_bottom_in[114], chany_bottom_in[155], chany_bottom_in[178]}),
		.sram(mux_tree_tapbuf_size8_43_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_43_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size8 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[77], chany_top_in[141], chany_bottom_in[46], chany_bottom_in[110], chany_bottom_in[143], chany_bottom_in[174]}),
		.sram(mux_tree_tapbuf_size8_44_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_44_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size8 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[78], chany_top_in[142], chany_bottom_in[45], chany_bottom_in[109], chany_bottom_in[139], chany_bottom_in[173]}),
		.sram(mux_tree_tapbuf_size8_45_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_45_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size8 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[80], chany_top_in[144], chany_bottom_in[44], chany_bottom_in[108], chany_bottom_in[135], chany_bottom_in[172]}),
		.sram(mux_tree_tapbuf_size8_46_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_46_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size8 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[81], chany_top_in[145], chany_bottom_in[42], chany_bottom_in[106], chany_bottom_in[131], chany_bottom_in[170]}),
		.sram(mux_tree_tapbuf_size8_47_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_47_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size8 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[82], chany_top_in[146], chany_bottom_in[41], chany_bottom_in[105], chany_bottom_in[127], chany_bottom_in[169]}),
		.sram(mux_tree_tapbuf_size8_48_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_48_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size8 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[84], chany_top_in[148], chany_bottom_in[40], chany_bottom_in[104], chany_bottom_in[123], chany_bottom_in[168]}),
		.sram(mux_tree_tapbuf_size8_49_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_49_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size8 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[85], chany_top_in[149], chany_bottom_in[38], chany_bottom_in[102], chany_bottom_in[119], chany_bottom_in[166]}),
		.sram(mux_tree_tapbuf_size8_50_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_50_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size8 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[89], chany_top_in[153], chany_bottom_in[34], chany_bottom_in[98], chany_bottom_in[107], chany_bottom_in[162]}),
		.sram(mux_tree_tapbuf_size8_51_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_51_sram_inv[0:3]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size8 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[90], chany_top_in[154], chany_bottom_in[33], chany_bottom_in[97], chany_bottom_in[103], chany_bottom_in[161]}),
		.sram(mux_tree_tapbuf_size8_52_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_52_sram_inv[0:3]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size8 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[92], chany_top_in[156], chany_bottom_in[32], chany_bottom_in[96], chany_bottom_in[99], chany_bottom_in[160]}),
		.sram(mux_tree_tapbuf_size8_53_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_53_sram_inv[0:3]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size8 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[93], chany_top_in[157], chany_bottom_in[30], chany_bottom_in[94:95], chany_bottom_in[158]}),
		.sram(mux_tree_tapbuf_size8_54_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_54_sram_inv[0:3]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size8 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[94:95], chany_top_in[158], chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[93], chany_bottom_in[157]}),
		.sram(mux_tree_tapbuf_size8_55_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_55_sram_inv[0:3]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size8 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[96], chany_top_in[99], chany_top_in[160], chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[92], chany_bottom_in[156]}),
		.sram(mux_tree_tapbuf_size8_56_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_56_sram_inv[0:3]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size8 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[97], chany_top_in[103], chany_top_in[161], chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[90], chany_bottom_in[154]}),
		.sram(mux_tree_tapbuf_size8_57_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_57_sram_inv[0:3]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size8 mux_right_track_232 (
		.in({chany_top_in[37], chany_top_in[101], chany_top_in[115], chany_top_in[165], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[86], chany_bottom_in[150]}),
		.sram(mux_tree_tapbuf_size8_58_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_58_sram_inv[0:3]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size8 mux_right_track_240 (
		.in({chany_top_in[38], chany_top_in[102], chany_top_in[119], chany_top_in[166], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[85], chany_bottom_in[149]}),
		.sram(mux_tree_tapbuf_size8_59_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_59_sram_inv[0:3]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size8 mux_right_track_248 (
		.in({chany_top_in[40], chany_top_in[104], chany_top_in[123], chany_top_in[168], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[84], chany_bottom_in[148]}),
		.sram(mux_tree_tapbuf_size8_60_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_60_sram_inv[0:3]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size8 mux_right_track_256 (
		.in({chany_top_in[41], chany_top_in[105], chany_top_in[127], chany_top_in[169], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[82], chany_bottom_in[146]}),
		.sram(mux_tree_tapbuf_size8_61_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_61_sram_inv[0:3]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size8 mux_right_track_264 (
		.in({chany_top_in[42], chany_top_in[106], chany_top_in[131], chany_top_in[170], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[81], chany_bottom_in[145]}),
		.sram(mux_tree_tapbuf_size8_62_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_62_sram_inv[0:3]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size8 mux_right_track_272 (
		.in({chany_top_in[44], chany_top_in[108], chany_top_in[135], chany_top_in[172], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[80], chany_bottom_in[144]}),
		.sram(mux_tree_tapbuf_size8_63_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_63_sram_inv[0:3]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size8 mux_right_track_280 (
		.in({chany_top_in[45], chany_top_in[109], chany_top_in[139], chany_top_in[173], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[78], chany_bottom_in[142]}),
		.sram(mux_tree_tapbuf_size8_64_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_64_sram_inv[0:3]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size8 mux_right_track_304 (
		.in({chany_top_in[49], chany_top_in[113], chany_top_in[151], chany_top_in[177], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[74], chany_bottom_in[138]}),
		.sram(mux_tree_tapbuf_size8_65_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_65_sram_inv[0:3]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size8 mux_right_track_312 (
		.in({chany_top_in[50], chany_top_in[114], chany_top_in[155], chany_top_in[178], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[73], chany_bottom_in[137]}),
		.sram(mux_tree_tapbuf_size8_66_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_66_sram_inv[0:3]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size8 mux_right_track_320 (
		.in({chany_top_in[52], chany_top_in[116], chany_top_in[159], chany_top_in[180], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[72], chany_bottom_in[136]}),
		.sram(mux_tree_tapbuf_size8_67_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_67_sram_inv[0:3]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size8 mux_right_track_328 (
		.in({chany_top_in[53], chany_top_in[117], chany_top_in[163], chany_top_in[181], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[70], chany_bottom_in[134]}),
		.sram(mux_tree_tapbuf_size8_68_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_68_sram_inv[0:3]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size8 mux_right_track_336 (
		.in({chany_top_in[54], chany_top_in[118], chany_top_in[167], chany_top_in[182], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[69], chany_bottom_in[133]}),
		.sram(mux_tree_tapbuf_size8_69_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_69_sram_inv[0:3]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size8 mux_right_track_344 (
		.in({chany_top_in[56], chany_top_in[120], chany_top_in[171], chany_top_in[184], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[68], chany_bottom_in[132]}),
		.sram(mux_tree_tapbuf_size8_70_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_70_sram_inv[0:3]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size8 mux_right_track_352 (
		.in({chany_top_in[57], chany_top_in[121], chany_top_in[175], chany_top_in[185], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[66], chany_bottom_in[130]}),
		.sram(mux_tree_tapbuf_size8_71_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_71_sram_inv[0:3]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size8 mux_right_track_368 (
		.in({chany_top_in[60], chany_top_in[124], chany_top_in[183], right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[64], chany_bottom_in[128]}),
		.sram(mux_tree_tapbuf_size8_72_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_72_sram_inv[0:3]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size8_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_0_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_1_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_2_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_3_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_4_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_5_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_6_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_7_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_8_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_9_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_10_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_11_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_12_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_13_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_14_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_15_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_16_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_17_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_18_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_19_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_20_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_21_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_22_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_23_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_24_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_25_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_26_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_27_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_28_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_29_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_30_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_31_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_32_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_33_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_34_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_35_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_36_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_37_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_38_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_39_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_39_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_40_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_40_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_41_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_41_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_42_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_42_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_43_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_43_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_44_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_44_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_45_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_45_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_46_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_46_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_47_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_47_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_48_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_48_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_49_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_49_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_50_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_50_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_51_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_51_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_52_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_52_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_53_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_53_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_54_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_54_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_55_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_55_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_56_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_56_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_57_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_57_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_58_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_58_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_59_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_59_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_60_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_60_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_61_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_61_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_62_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_62_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_63_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_63_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_64_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_64_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_65_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_65_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_66_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_66_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_67_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_67_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_68_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_68_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_69_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_69_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_70_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_70_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_71_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_71_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_72_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_72_sram_inv[0:3]));

	mux_tree_tapbuf_size7 mux_top_track_16 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[68], chanx_right_in[132], chanx_left_in[61], chanx_left_in[125], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size7 mux_top_track_24 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[69], chanx_right_in[133], chanx_left_in[60], chanx_left_in[124], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size7 mux_top_track_352 (
		.in({chanx_right_in[60], chanx_right_in[124], chanx_right_in[183], chanx_left_in[5], chanx_left_in[19], chanx_left_in[69], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size7 mux_right_track_0 (
		.in({chany_top_in[62], chany_top_in[126], chany_top_in[188], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, chany_bottom_in[61], chany_bottom_in[125], chany_bottom_in[187]}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size7_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_right_track_376 (
		.in({chany_top_in[61], chany_top_in[125], chany_top_in[187], chany_bottom_in[62], chany_bottom_in[126], chany_bottom_in[188]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size6_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size19 mux_bottom_track_1 (
		.in({chanx_right_in[61], chanx_right_in[125], chanx_right_in[187], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[1], chanx_left_in[7], chanx_left_in[65], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size19_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_0_sram_inv[0:4]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size19 mux_bottom_track_9 (
		.in({chanx_right_in[60], chanx_right_in[124], chanx_right_in[183], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[2], chanx_left_in[11], chanx_left_in[66], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size19_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_1_sram_inv[0:4]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size19 mux_bottom_track_17 (
		.in({chanx_right_in[58], chanx_right_in[122], chanx_right_in[179], chanx_right_in[186], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[4], chanx_left_in[15], chanx_left_in[68], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size19_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_2_sram_inv[0:4]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size19 mux_bottom_track_25 (
		.in({chanx_right_in[57], chanx_right_in[121], chanx_right_in[175], chanx_right_in[185], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[5], chanx_left_in[19], chanx_left_in[69], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size19_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_3_sram_inv[0:4]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size19 mux_bottom_track_33 (
		.in({chanx_right_in[56], chanx_right_in[120], chanx_right_in[171], chanx_right_in[184], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[6], chanx_left_in[23], chanx_left_in[70], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size19_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_4_sram_inv[0:4]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size19 mux_bottom_track_41 (
		.in({chanx_right_in[54], chanx_right_in[118], chanx_right_in[167], chanx_right_in[182], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[8], chanx_left_in[27], chanx_left_in[72], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size19_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_5_sram_inv[0:4]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size19 mux_bottom_track_49 (
		.in({chanx_right_in[53], chanx_right_in[117], chanx_right_in[163], chanx_right_in[181], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[9], chanx_left_in[31], chanx_left_in[73], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size19_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_6_sram_inv[0:4]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size19 mux_bottom_track_57 (
		.in({chanx_right_in[52], chanx_right_in[116], chanx_right_in[159], chanx_right_in[180], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[10], chanx_left_in[35], chanx_left_in[74], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size19_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_7_sram_inv[0:4]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size19 mux_bottom_track_65 (
		.in({chanx_right_in[50], chanx_right_in[114], chanx_right_in[155], chanx_right_in[178], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[12], chanx_left_in[39], chanx_left_in[76], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size19_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_8_sram_inv[0:4]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size19 mux_bottom_track_89 (
		.in({chanx_right_in[46], chanx_right_in[110], chanx_right_in[143], chanx_right_in[174], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[16], chanx_left_in[51], chanx_left_in[80], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size19_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_9_sram_inv[0:4]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size19 mux_bottom_track_97 (
		.in({chanx_right_in[45], chanx_right_in[109], chanx_right_in[139], chanx_right_in[173], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[17], chanx_left_in[55], chanx_left_in[81], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size19_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_10_sram_inv[0:4]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size19 mux_bottom_track_105 (
		.in({chanx_right_in[44], chanx_right_in[108], chanx_right_in[135], chanx_right_in[172], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[18], chanx_left_in[59], chanx_left_in[82], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size19_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_11_sram_inv[0:4]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size19 mux_bottom_track_113 (
		.in({chanx_right_in[42], chanx_right_in[106], chanx_right_in[131], chanx_right_in[170], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[20], chanx_left_in[63], chanx_left_in[84], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size19_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_12_sram_inv[0:4]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size19 mux_bottom_track_121 (
		.in({chanx_right_in[41], chanx_right_in[105], chanx_right_in[127], chanx_right_in[169], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[21], chanx_left_in[67], chanx_left_in[85], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size19_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_13_sram_inv[0:4]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size19 mux_bottom_track_129 (
		.in({chanx_right_in[40], chanx_right_in[104], chanx_right_in[123], chanx_right_in[168], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[22], chanx_left_in[71], chanx_left_in[86], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size19_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_14_sram_inv[0:4]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size19 mux_bottom_track_137 (
		.in({chanx_right_in[38], chanx_right_in[102], chanx_right_in[119], chanx_right_in[166], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[24], chanx_left_in[75], chanx_left_in[88], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size19_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_15_sram_inv[0:4]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size19 mux_bottom_track_161 (
		.in({chanx_right_in[34], chanx_right_in[98], chanx_right_in[107], chanx_right_in[162], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[28], chanx_left_in[87], chanx_left_in[92], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size19_16_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_16_sram_inv[0:4]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size19 mux_bottom_track_169 (
		.in({chanx_right_in[33], chanx_right_in[97], chanx_right_in[103], chanx_right_in[161], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[29], chanx_left_in[91], chanx_left_in[93], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size19_17_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_17_sram_inv[0:4]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size19 mux_bottom_track_177 (
		.in({chanx_right_in[32], chanx_right_in[96], chanx_right_in[99], chanx_right_in[160], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[30], chanx_left_in[94:95], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size19_18_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_18_sram_inv[0:4]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size19 mux_bottom_track_185 (
		.in({chanx_right_in[30], chanx_right_in[94:95], chanx_right_in[158], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[32], chanx_left_in[96], chanx_left_in[99], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size19_19_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_19_sram_inv[0:4]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size19 mux_bottom_track_193 (
		.in({chanx_right_in[29], chanx_right_in[91], chanx_right_in[93], chanx_right_in[157], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[33], chanx_left_in[97], chanx_left_in[103], chanx_left_in[161]}),
		.sram(mux_tree_tapbuf_size19_20_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_20_sram_inv[0:4]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size19 mux_bottom_track_201 (
		.in({chanx_right_in[28], chanx_right_in[87], chanx_right_in[92], chanx_right_in[156], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[34], chanx_left_in[98], chanx_left_in[107], chanx_left_in[162]}),
		.sram(mux_tree_tapbuf_size19_21_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_21_sram_inv[0:4]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size19 mux_bottom_track_209 (
		.in({chanx_right_in[26], chanx_right_in[83], chanx_right_in[90], chanx_right_in[154], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[36], chanx_left_in[100], chanx_left_in[111], chanx_left_in[164]}),
		.sram(mux_tree_tapbuf_size19_22_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_22_sram_inv[0:4]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size19 mux_bottom_track_233 (
		.in({chanx_right_in[22], chanx_right_in[71], chanx_right_in[86], chanx_right_in[150], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[40], chanx_left_in[104], chanx_left_in[123], chanx_left_in[168]}),
		.sram(mux_tree_tapbuf_size19_23_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_23_sram_inv[0:4]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size19 mux_bottom_track_241 (
		.in({chanx_right_in[21], chanx_right_in[67], chanx_right_in[85], chanx_right_in[149], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[41], chanx_left_in[105], chanx_left_in[127], chanx_left_in[169]}),
		.sram(mux_tree_tapbuf_size19_24_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_24_sram_inv[0:4]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size19 mux_bottom_track_249 (
		.in({chanx_right_in[20], chanx_right_in[63], chanx_right_in[84], chanx_right_in[148], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[42], chanx_left_in[106], chanx_left_in[131], chanx_left_in[170]}),
		.sram(mux_tree_tapbuf_size19_25_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_25_sram_inv[0:4]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size19 mux_bottom_track_257 (
		.in({chanx_right_in[18], chanx_right_in[59], chanx_right_in[82], chanx_right_in[146], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[44], chanx_left_in[108], chanx_left_in[135], chanx_left_in[172]}),
		.sram(mux_tree_tapbuf_size19_26_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_26_sram_inv[0:4]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size19 mux_bottom_track_265 (
		.in({chanx_right_in[17], chanx_right_in[55], chanx_right_in[81], chanx_right_in[145], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[45], chanx_left_in[109], chanx_left_in[139], chanx_left_in[173]}),
		.sram(mux_tree_tapbuf_size19_27_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_27_sram_inv[0:4]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size19 mux_bottom_track_273 (
		.in({chanx_right_in[16], chanx_right_in[51], chanx_right_in[80], chanx_right_in[144], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[46], chanx_left_in[110], chanx_left_in[143], chanx_left_in[174]}),
		.sram(mux_tree_tapbuf_size19_28_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_28_sram_inv[0:4]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size19 mux_bottom_track_281 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[78], chanx_right_in[142], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[48], chanx_left_in[112], chanx_left_in[147], chanx_left_in[176]}),
		.sram(mux_tree_tapbuf_size19_29_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_29_sram_inv[0:4]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size19 mux_bottom_track_305 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[74], chanx_right_in[138], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[52], chanx_left_in[116], chanx_left_in[159], chanx_left_in[180]}),
		.sram(mux_tree_tapbuf_size19_30_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_30_sram_inv[0:4]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size19 mux_bottom_track_313 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[73], chanx_right_in[137], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_7_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_199_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[53], chanx_left_in[117], chanx_left_in[163], chanx_left_in[181]}),
		.sram(mux_tree_tapbuf_size19_31_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_31_sram_inv[0:4]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size19 mux_bottom_track_321 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[72], chanx_right_in[136], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_11_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_203_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[54], chanx_left_in[118], chanx_left_in[167], chanx_left_in[182]}),
		.sram(mux_tree_tapbuf_size19_32_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_32_sram_inv[0:4]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size19 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[64], chany_top_in[128], chany_bottom_in[62], chany_bottom_in[126], chany_bottom_in[188], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size19_33_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_33_sram_inv[0:4]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size19 mux_left_track_33 (
		.in({chany_top_in[58], chany_top_in[122], chany_top_in[179], chany_top_in[186], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[68], chany_bottom_in[132], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size19_34_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_34_sram_inv[0:4]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size19 mux_left_track_41 (
		.in({chany_top_in[57], chany_top_in[121], chany_top_in[175], chany_top_in[185], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[69], chany_bottom_in[133], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size19_35_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_35_sram_inv[0:4]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size19 mux_left_track_49 (
		.in({chany_top_in[56], chany_top_in[120], chany_top_in[171], chany_top_in[184], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[70], chany_bottom_in[134], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size19_36_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_36_sram_inv[0:4]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size19 mux_left_track_57 (
		.in({chany_top_in[54], chany_top_in[118], chany_top_in[167], chany_top_in[182], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[72], chany_bottom_in[136], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size19_37_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_37_sram_inv[0:4]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size19 mux_left_track_65 (
		.in({chany_top_in[53], chany_top_in[117], chany_top_in[163], chany_top_in[181], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[73], chany_bottom_in[137], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size19_38_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_38_sram_inv[0:4]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size19 mux_left_track_81 (
		.in({chany_top_in[50], chany_top_in[114], chany_top_in[155], chany_top_in[178], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[76], chany_bottom_in[140], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size19_39_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_39_sram_inv[0:4]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size19 mux_left_track_89 (
		.in({chany_top_in[49], chany_top_in[113], chany_top_in[151], chany_top_in[177], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[77], chany_bottom_in[141], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size19_40_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_40_sram_inv[0:4]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size19 mux_left_track_97 (
		.in({chany_top_in[48], chany_top_in[112], chany_top_in[147], chany_top_in[176], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[78], chany_bottom_in[142], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size19_41_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_41_sram_inv[0:4]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size19 mux_left_track_105 (
		.in({chany_top_in[46], chany_top_in[110], chany_top_in[143], chany_top_in[174], chany_bottom_in[16], chany_bottom_in[51], chany_bottom_in[80], chany_bottom_in[144], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size19_42_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_42_sram_inv[0:4]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size19 mux_left_track_113 (
		.in({chany_top_in[45], chany_top_in[109], chany_top_in[139], chany_top_in[173], chany_bottom_in[17], chany_bottom_in[55], chany_bottom_in[81], chany_bottom_in[145], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size19_43_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_43_sram_inv[0:4]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size19 mux_left_track_121 (
		.in({chany_top_in[44], chany_top_in[108], chany_top_in[135], chany_top_in[172], chany_bottom_in[18], chany_bottom_in[59], chany_bottom_in[82], chany_bottom_in[146], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size19_44_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_44_sram_inv[0:4]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size19 mux_left_track_129 (
		.in({chany_top_in[42], chany_top_in[106], chany_top_in[131], chany_top_in[170], chany_bottom_in[20], chany_bottom_in[63], chany_bottom_in[84], chany_bottom_in[148], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size19_45_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_45_sram_inv[0:4]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size19 mux_left_track_137 (
		.in({chany_top_in[41], chany_top_in[105], chany_top_in[127], chany_top_in[169], chany_bottom_in[21], chany_bottom_in[67], chany_bottom_in[85], chany_bottom_in[149], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size19_46_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_46_sram_inv[0:4]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size19 mux_left_track_153 (
		.in({chany_top_in[38], chany_top_in[102], chany_top_in[119], chany_top_in[166], chany_bottom_in[24], chany_bottom_in[75], chany_bottom_in[88], chany_bottom_in[152], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size19_47_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_47_sram_inv[0:4]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size19 mux_left_track_161 (
		.in({chany_top_in[37], chany_top_in[101], chany_top_in[115], chany_top_in[165], chany_bottom_in[25], chany_bottom_in[79], chany_bottom_in[89], chany_bottom_in[153], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size19_48_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_48_sram_inv[0:4]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size19 mux_left_track_169 (
		.in({chany_top_in[36], chany_top_in[100], chany_top_in[111], chany_top_in[164], chany_bottom_in[26], chany_bottom_in[83], chany_bottom_in[90], chany_bottom_in[154], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size19_49_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_49_sram_inv[0:4]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size19 mux_left_track_177 (
		.in({chany_top_in[34], chany_top_in[98], chany_top_in[107], chany_top_in[162], chany_bottom_in[28], chany_bottom_in[87], chany_bottom_in[92], chany_bottom_in[156], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size19_50_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_50_sram_inv[0:4]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size19 mux_left_track_185 (
		.in({chany_top_in[33], chany_top_in[97], chany_top_in[103], chany_top_in[161], chany_bottom_in[29], chany_bottom_in[91], chany_bottom_in[93], chany_bottom_in[157], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size19_51_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_51_sram_inv[0:4]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size19 mux_left_track_193 (
		.in({chany_top_in[32], chany_top_in[96], chany_top_in[99], chany_top_in[160], chany_bottom_in[30], chany_bottom_in[94:95], chany_bottom_in[158], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size19_52_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_52_sram_inv[0:4]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size19 mux_left_track_201 (
		.in({chany_top_in[30], chany_top_in[94:95], chany_top_in[158], chany_bottom_in[32], chany_bottom_in[96], chany_bottom_in[99], chany_bottom_in[160], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size19_53_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_53_sram_inv[0:4]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size19 mux_left_track_209 (
		.in({chany_top_in[29], chany_top_in[91], chany_top_in[93], chany_top_in[157], chany_bottom_in[33], chany_bottom_in[97], chany_bottom_in[103], chany_bottom_in[161], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size19_54_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_54_sram_inv[0:4]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size19 mux_left_track_225 (
		.in({chany_top_in[26], chany_top_in[83], chany_top_in[90], chany_top_in[154], chany_bottom_in[36], chany_bottom_in[100], chany_bottom_in[111], chany_bottom_in[164], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size19_55_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_55_sram_inv[0:4]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size19 mux_left_track_233 (
		.in({chany_top_in[25], chany_top_in[79], chany_top_in[89], chany_top_in[153], chany_bottom_in[37], chany_bottom_in[101], chany_bottom_in[115], chany_bottom_in[165], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size19_56_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_56_sram_inv[0:4]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size19 mux_left_track_241 (
		.in({chany_top_in[24], chany_top_in[75], chany_top_in[88], chany_top_in[152], chany_bottom_in[38], chany_bottom_in[102], chany_bottom_in[119], chany_bottom_in[166], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size19_57_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_57_sram_inv[0:4]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size19 mux_left_track_249 (
		.in({chany_top_in[22], chany_top_in[71], chany_top_in[86], chany_top_in[150], chany_bottom_in[40], chany_bottom_in[104], chany_bottom_in[123], chany_bottom_in[168], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size19_58_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_58_sram_inv[0:4]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size19 mux_left_track_257 (
		.in({chany_top_in[21], chany_top_in[67], chany_top_in[85], chany_top_in[149], chany_bottom_in[41], chany_bottom_in[105], chany_bottom_in[127], chany_bottom_in[169], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size19_59_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_59_sram_inv[0:4]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size19 mux_left_track_265 (
		.in({chany_top_in[20], chany_top_in[63], chany_top_in[84], chany_top_in[148], chany_bottom_in[42], chany_bottom_in[106], chany_bottom_in[131], chany_bottom_in[170], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size19_60_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_60_sram_inv[0:4]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size19 mux_left_track_273 (
		.in({chany_top_in[18], chany_top_in[59], chany_top_in[82], chany_top_in[146], chany_bottom_in[44], chany_bottom_in[108], chany_bottom_in[135], chany_bottom_in[172], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size19_61_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_61_sram_inv[0:4]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size19 mux_left_track_281 (
		.in({chany_top_in[17], chany_top_in[55], chany_top_in[81], chany_top_in[145], chany_bottom_in[45], chany_bottom_in[109], chany_bottom_in[139], chany_bottom_in[173], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size19_62_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_62_sram_inv[0:4]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size19 mux_left_track_297 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[78], chany_top_in[142], chany_bottom_in[48], chany_bottom_in[112], chany_bottom_in[147], chany_bottom_in[176], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size19_63_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_63_sram_inv[0:4]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size19 mux_left_track_305 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[77], chany_top_in[141], chany_bottom_in[49], chany_bottom_in[113], chany_bottom_in[151], chany_bottom_in[177], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size19_64_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_64_sram_inv[0:4]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size19 mux_left_track_313 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[76], chany_top_in[140], chany_bottom_in[50], chany_bottom_in[114], chany_bottom_in[155], chany_bottom_in[178], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size19_65_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_65_sram_inv[0:4]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size19 mux_left_track_361 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[68], chany_top_in[132], chany_bottom_in[58], chany_bottom_in[122], chany_bottom_in[179], chany_bottom_in[186], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size19_66_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size19_66_sram_inv[0:4]),
		.out(chanx_left_out[180]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_0_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_1_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_2_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_3_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_4_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_5_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_6_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_7_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_8_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_9_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_10_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_11_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_12_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_13_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_14_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_15_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_16_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_16_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_17_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_17_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_18_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_18_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_19_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_19_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_20_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_20_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_21_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_21_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_22_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_22_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_23_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_23_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_24_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_24_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_25_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_25_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_26_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_26_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_27_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_27_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_28_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_28_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_29_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_29_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_30_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_30_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_31_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_31_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_32_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_32_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_33_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_33_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_34_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_34_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_35_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_35_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_36_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_36_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_37_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_37_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_38_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_38_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_39_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_39_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_40_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_40_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_41_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_41_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_42_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_42_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_43_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_43_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_44_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_44_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_45_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_45_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_46_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_46_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_47_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_47_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_48_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_48_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_49_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_49_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_50_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_50_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_51_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_51_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_52_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_52_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_53_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_53_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_54_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_54_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_55_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_55_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_56_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_56_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_57_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_57_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_58_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_58_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_59_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_59_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_60_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_60_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_61_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_61_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_62_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_62_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_63_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_63_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_64_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_64_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_65_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_65_sram_inv[0:4]));

	mux_tree_tapbuf_size19_mem mem_left_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size19_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size19_66_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size19_66_sram_inv[0:4]));

	mux_tree_tapbuf_size20 mux_bottom_track_73 (
		.in({chanx_right_in[49], chanx_right_in[113], chanx_right_in[151], chanx_right_in[177], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_43_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_235_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[13], chanx_left_in[43], chanx_left_in[77], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size20_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_0_sram_inv[0:4]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size20 mux_bottom_track_81 (
		.in({chanx_right_in[48], chanx_right_in[112], chanx_right_in[147], chanx_right_in[176], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_47_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_239_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[14], chanx_left_in[47], chanx_left_in[78], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size20_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_1_sram_inv[0:4]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size20 mux_bottom_track_145 (
		.in({chanx_right_in[37], chanx_right_in[101], chanx_right_in[115], chanx_right_in[165], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_79_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_271_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[25], chanx_left_in[79], chanx_left_in[89], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size20_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_2_sram_inv[0:4]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size20 mux_bottom_track_153 (
		.in({chanx_right_in[36], chanx_right_in[100], chanx_right_in[111], chanx_right_in[164], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_83_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_275_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[26], chanx_left_in[83], chanx_left_in[90], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size20_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_3_sram_inv[0:4]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size20 mux_bottom_track_217 (
		.in({chanx_right_in[25], chanx_right_in[79], chanx_right_in[89], chanx_right_in[153], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_115_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_307_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[37], chanx_left_in[101], chanx_left_in[115], chanx_left_in[165]}),
		.sram(mux_tree_tapbuf_size20_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_4_sram_inv[0:4]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size20 mux_bottom_track_225 (
		.in({chanx_right_in[24], chanx_right_in[75], chanx_right_in[88], chanx_right_in[152], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_119_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_311_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[38], chanx_left_in[102], chanx_left_in[119], chanx_left_in[166]}),
		.sram(mux_tree_tapbuf_size20_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_5_sram_inv[0:4]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size20 mux_bottom_track_289 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[77], chanx_right_in[141], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_151_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_3_, chanx_left_in[49], chanx_left_in[113], chanx_left_in[151], chanx_left_in[177]}),
		.sram(mux_tree_tapbuf_size20_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_6_sram_inv[0:4]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size20 mux_bottom_track_297 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[76], chanx_right_in[140], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_155_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_7_, chanx_left_in[50], chanx_left_in[114], chanx_left_in[155], chanx_left_in[178]}),
		.sram(mux_tree_tapbuf_size20_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_7_sram_inv[0:4]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size20 mux_left_track_73 (
		.in({chany_top_in[52], chany_top_in[116], chany_top_in[159], chany_top_in[180], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[74], chany_bottom_in[138], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size20_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_8_sram_inv[0:4]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size20 mux_left_track_145 (
		.in({chany_top_in[40], chany_top_in[104], chany_top_in[123], chany_top_in[168], chany_bottom_in[22], chany_bottom_in[71], chany_bottom_in[86], chany_bottom_in[150], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size20_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_9_sram_inv[0:4]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size20 mux_left_track_217 (
		.in({chany_top_in[28], chany_top_in[87], chany_top_in[92], chany_top_in[156], chany_bottom_in[34], chany_bottom_in[98], chany_bottom_in[107], chany_bottom_in[162], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size20_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_10_sram_inv[0:4]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size20 mux_left_track_289 (
		.in({chany_top_in[16], chany_top_in[51], chany_top_in[80], chany_top_in[144], chany_bottom_in[46], chany_bottom_in[110], chany_bottom_in[143], chany_bottom_in[174], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size20_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_11_sram_inv[0:4]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_0_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_1_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_2_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_3_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_4_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_5_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_6_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_7_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_8_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_9_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_10_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_11_sram_inv[0:4]));

	mux_tree_tapbuf_size18 mux_bottom_track_329 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[70], chanx_right_in[134], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_15_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_51_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_87_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_123_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_159_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_207_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_243_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_279_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_315_, chanx_left_in[56], chanx_left_in[120], chanx_left_in[171], chanx_left_in[184]}),
		.sram(mux_tree_tapbuf_size18_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_0_sram_inv[0:4]),
		.out(chany_bottom_out[164]));

	mux_tree_tapbuf_size18 mux_bottom_track_337 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[69], chanx_right_in[133], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_19_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_55_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_91_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_127_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_163_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_211_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_247_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_283_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_319_, chanx_left_in[57], chanx_left_in[121], chanx_left_in[175], chanx_left_in[185]}),
		.sram(mux_tree_tapbuf_size18_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_1_sram_inv[0:4]),
		.out(chany_bottom_out[168]));

	mux_tree_tapbuf_size18 mux_bottom_track_345 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[68], chanx_right_in[132], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_23_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_59_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_95_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_131_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_167_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_215_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_251_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_287_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_323_, chanx_left_in[58], chanx_left_in[122], chanx_left_in[179], chanx_left_in[186]}),
		.sram(mux_tree_tapbuf_size18_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_2_sram_inv[0:4]),
		.out(chany_bottom_out[172]));

	mux_tree_tapbuf_size18 mux_bottom_track_361 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[65], chanx_right_in[129], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_31_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_67_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_103_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_139_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_175_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_187_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_223_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_259_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_295_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_331_, chanx_left_in[61], chanx_left_in[125], chanx_left_in[187]}),
		.sram(mux_tree_tapbuf_size18_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_3_sram_inv[0:4]),
		.out(chany_bottom_out[180]));

	mux_tree_tapbuf_size18 mux_bottom_track_369 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[64], chanx_right_in[128], bottom_left_grid_right_width_0_height_0_subtile_0__pin_error_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_35_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_71_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_107_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_143_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_179_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_191_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_227_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_263_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_299_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_335_, chanx_left_in[62], chanx_left_in[126], chanx_left_in[188]}),
		.sram(mux_tree_tapbuf_size18_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_4_sram_inv[0:4]),
		.out(chany_bottom_out[184]));

	mux_tree_tapbuf_size18 mux_bottom_track_377 (
		.in({chanx_right_in[62], chanx_right_in[126], chanx_right_in[188], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_3_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_39_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_75_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_111_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_147_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_195_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_231_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_267_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_303_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_339_, chanx_left_in[0], chanx_left_in[3], chanx_left_in[64], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size18_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_5_sram_inv[0:4]),
		.out(chany_bottom_out[188]));

	mux_tree_tapbuf_size18 mux_left_track_9 (
		.in({chany_top_in[62], chany_top_in[126], chany_top_in[188], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[64], chany_bottom_in[128], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size18_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_6_sram_inv[0:4]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size18 mux_left_track_17 (
		.in({chany_top_in[61], chany_top_in[125], chany_top_in[187], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[65], chany_bottom_in[129], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size18_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_7_sram_inv[0:4]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size18 mux_left_track_25 (
		.in({chany_top_in[60], chany_top_in[124], chany_top_in[183], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[66], chany_bottom_in[130], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size18_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_8_sram_inv[0:4]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size18 mux_left_track_321 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[74], chany_top_in[138], chany_bottom_in[52], chany_bottom_in[116], chany_bottom_in[159], chany_bottom_in[180], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size18_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_9_sram_inv[0:4]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size18 mux_left_track_329 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[73], chany_top_in[137], chany_bottom_in[53], chany_bottom_in[117], chany_bottom_in[163], chany_bottom_in[181], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size18_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_10_sram_inv[0:4]),
		.out(chanx_left_out[164]));

	mux_tree_tapbuf_size18 mux_left_track_337 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[72], chany_top_in[136], chany_bottom_in[54], chany_bottom_in[118], chany_bottom_in[167], chany_bottom_in[182], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size18_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_11_sram_inv[0:4]),
		.out(chanx_left_out[168]));

	mux_tree_tapbuf_size18 mux_left_track_345 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[70], chany_top_in[134], chany_bottom_in[56], chany_bottom_in[120], chany_bottom_in[171], chany_bottom_in[184], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size18_12_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_12_sram_inv[0:4]),
		.out(chanx_left_out[172]));

	mux_tree_tapbuf_size18 mux_left_track_353 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[69], chany_top_in[133], chany_bottom_in[57], chany_bottom_in[121], chany_bottom_in[175], chany_bottom_in[185], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size18_13_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_13_sram_inv[0:4]),
		.out(chanx_left_out[176]));

	mux_tree_tapbuf_size18 mux_left_track_369 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[66], chany_top_in[130], chany_bottom_in[60], chany_bottom_in[124], chany_bottom_in[183], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size18_14_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_14_sram_inv[0:4]),
		.out(chanx_left_out[184]));

	mux_tree_tapbuf_size18 mux_left_track_377 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[65], chany_top_in[129], chany_bottom_in[61], chany_bottom_in[125], chany_bottom_in[187], left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size18_15_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size18_15_sram_inv[0:4]),
		.out(chanx_left_out[188]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_0_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_1_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_2_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_361 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_3_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_4_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_bottom_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_5_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_6_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_7_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_8_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_9_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_329 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_10_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_337 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_11_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_345 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_12_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_12_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_13_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_13_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_369 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size19_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size18_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_14_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_14_sram_inv[0:4]));

	mux_tree_tapbuf_size18_mem mem_left_track_377 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_14_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size18_15_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size18_15_sram_inv[0:4]));

	mux_tree_tapbuf_size17 mux_bottom_track_353 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[66], chanx_right_in[130], bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_27_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_63_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_99_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_135_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_171_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_183_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_219_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_255_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_291_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_channel_out_op_327_, chanx_left_in[60], chanx_left_in[124], chanx_left_in[183]}),
		.sram(mux_tree_tapbuf_size17_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size17_0_sram_inv[0:4]),
		.out(chany_bottom_out[176]));

	mux_tree_tapbuf_size17_mem mem_bottom_track_353 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size18_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size17_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size17_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size17_0_sram_inv[0:4]));

endmodule
// ----- END Verilog module for sb_1__2_ -----

//----- Default net type -----
`default_nettype wire



