//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[5][5]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Wed Jul 24 20:28:26 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_5__5_ -----
module sb_5__5_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                chanx_left_in,
                left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                chanx_left_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:104] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_;
//----- INPUT PORTS -----
input [0:104] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:104] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:104] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:104] chany_top_out;
//----- OUTPUT PORTS -----
output [0:104] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:104] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:104] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_10_sram;
wire [0:3] mux_tree_tapbuf_size14_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_11_sram;
wire [0:3] mux_tree_tapbuf_size14_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_12_sram;
wire [0:3] mux_tree_tapbuf_size14_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_13_sram;
wire [0:3] mux_tree_tapbuf_size14_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_14_sram;
wire [0:3] mux_tree_tapbuf_size14_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_15_sram;
wire [0:3] mux_tree_tapbuf_size14_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_16_sram;
wire [0:3] mux_tree_tapbuf_size14_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_17_sram;
wire [0:3] mux_tree_tapbuf_size14_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_18_sram;
wire [0:3] mux_tree_tapbuf_size14_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_19_sram;
wire [0:3] mux_tree_tapbuf_size14_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_1_sram;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_20_sram;
wire [0:3] mux_tree_tapbuf_size14_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_21_sram;
wire [0:3] mux_tree_tapbuf_size14_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_22_sram;
wire [0:3] mux_tree_tapbuf_size14_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_23_sram;
wire [0:3] mux_tree_tapbuf_size14_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_24_sram;
wire [0:3] mux_tree_tapbuf_size14_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_25_sram;
wire [0:3] mux_tree_tapbuf_size14_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_26_sram;
wire [0:3] mux_tree_tapbuf_size14_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_27_sram;
wire [0:3] mux_tree_tapbuf_size14_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_28_sram;
wire [0:3] mux_tree_tapbuf_size14_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_29_sram;
wire [0:3] mux_tree_tapbuf_size14_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_2_sram;
wire [0:3] mux_tree_tapbuf_size14_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_30_sram;
wire [0:3] mux_tree_tapbuf_size14_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_31_sram;
wire [0:3] mux_tree_tapbuf_size14_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_32_sram;
wire [0:3] mux_tree_tapbuf_size14_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_33_sram;
wire [0:3] mux_tree_tapbuf_size14_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_34_sram;
wire [0:3] mux_tree_tapbuf_size14_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_35_sram;
wire [0:3] mux_tree_tapbuf_size14_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_36_sram;
wire [0:3] mux_tree_tapbuf_size14_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_37_sram;
wire [0:3] mux_tree_tapbuf_size14_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_38_sram;
wire [0:3] mux_tree_tapbuf_size14_38_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_3_sram;
wire [0:3] mux_tree_tapbuf_size14_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_4_sram;
wire [0:3] mux_tree_tapbuf_size14_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_5_sram;
wire [0:3] mux_tree_tapbuf_size14_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_6_sram;
wire [0:3] mux_tree_tapbuf_size14_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_7_sram;
wire [0:3] mux_tree_tapbuf_size14_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_8_sram;
wire [0:3] mux_tree_tapbuf_size14_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_9_sram;
wire [0:3] mux_tree_tapbuf_size14_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size15_0_sram;
wire [0:3] mux_tree_tapbuf_size15_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_1_sram;
wire [0:3] mux_tree_tapbuf_size15_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_2_sram;
wire [0:3] mux_tree_tapbuf_size15_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_3_sram;
wire [0:3] mux_tree_tapbuf_size15_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size15_4_sram;
wire [0:3] mux_tree_tapbuf_size15_4_sram_inv;
wire [0:0] mux_tree_tapbuf_size15_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size15_mem_4_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_4_sram;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_5_sram;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_6_sram;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_7_sram;
wire [0:2] mux_tree_tapbuf_size7_7_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail;
wire [0:3] mux_tree_tapbuf_size8_0_sram;
wire [0:3] mux_tree_tapbuf_size8_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_10_sram;
wire [0:3] mux_tree_tapbuf_size8_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_11_sram;
wire [0:3] mux_tree_tapbuf_size8_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_12_sram;
wire [0:3] mux_tree_tapbuf_size8_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_13_sram;
wire [0:3] mux_tree_tapbuf_size8_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_14_sram;
wire [0:3] mux_tree_tapbuf_size8_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_15_sram;
wire [0:3] mux_tree_tapbuf_size8_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_16_sram;
wire [0:3] mux_tree_tapbuf_size8_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_17_sram;
wire [0:3] mux_tree_tapbuf_size8_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_18_sram;
wire [0:3] mux_tree_tapbuf_size8_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_19_sram;
wire [0:3] mux_tree_tapbuf_size8_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_1_sram;
wire [0:3] mux_tree_tapbuf_size8_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_20_sram;
wire [0:3] mux_tree_tapbuf_size8_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_21_sram;
wire [0:3] mux_tree_tapbuf_size8_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_22_sram;
wire [0:3] mux_tree_tapbuf_size8_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_23_sram;
wire [0:3] mux_tree_tapbuf_size8_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_24_sram;
wire [0:3] mux_tree_tapbuf_size8_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_25_sram;
wire [0:3] mux_tree_tapbuf_size8_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_26_sram;
wire [0:3] mux_tree_tapbuf_size8_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_27_sram;
wire [0:3] mux_tree_tapbuf_size8_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_28_sram;
wire [0:3] mux_tree_tapbuf_size8_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_29_sram;
wire [0:3] mux_tree_tapbuf_size8_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_2_sram;
wire [0:3] mux_tree_tapbuf_size8_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_30_sram;
wire [0:3] mux_tree_tapbuf_size8_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_31_sram;
wire [0:3] mux_tree_tapbuf_size8_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_32_sram;
wire [0:3] mux_tree_tapbuf_size8_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_33_sram;
wire [0:3] mux_tree_tapbuf_size8_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_34_sram;
wire [0:3] mux_tree_tapbuf_size8_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_35_sram;
wire [0:3] mux_tree_tapbuf_size8_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_36_sram;
wire [0:3] mux_tree_tapbuf_size8_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_37_sram;
wire [0:3] mux_tree_tapbuf_size8_37_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_3_sram;
wire [0:3] mux_tree_tapbuf_size8_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_4_sram;
wire [0:3] mux_tree_tapbuf_size8_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_5_sram;
wire [0:3] mux_tree_tapbuf_size8_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_6_sram;
wire [0:3] mux_tree_tapbuf_size8_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_7_sram;
wire [0:3] mux_tree_tapbuf_size8_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_8_sram;
wire [0:3] mux_tree_tapbuf_size8_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size8_9_sram;
wire [0:3] mux_tree_tapbuf_size8_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size8_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size8_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_1_sram;
wire [0:3] mux_tree_tapbuf_size9_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_2_sram;
wire [0:3] mux_tree_tapbuf_size9_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_3_sram;
wire [0:3] mux_tree_tapbuf_size9_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_4_sram;
wire [0:3] mux_tree_tapbuf_size9_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_5_sram;
wire [0:3] mux_tree_tapbuf_size9_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_6_sram;
wire [0:3] mux_tree_tapbuf_size9_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size9_7_sram;
wire [0:3] mux_tree_tapbuf_size9_7_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size9_mem_7_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 160 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[1] = chanx_right_in[0];
// ----- Local connection due to Wire 161 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[2] = chanx_right_in[1];
// ----- Local connection due to Wire 162 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[3] = chanx_right_in[2];
// ----- Local connection due to Wire 164 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[5] = chanx_right_in[4];
// ----- Local connection due to Wire 165 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[6] = chanx_right_in[5];
// ----- Local connection due to Wire 166 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[7] = chanx_right_in[6];
// ----- Local connection due to Wire 168 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[9] = chanx_right_in[8];
// ----- Local connection due to Wire 169 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[10] = chanx_right_in[9];
// ----- Local connection due to Wire 170 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[11] = chanx_right_in[10];
// ----- Local connection due to Wire 172 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[13] = chanx_right_in[12];
// ----- Local connection due to Wire 173 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[14] = chanx_right_in[13];
// ----- Local connection due to Wire 174 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[15] = chanx_right_in[14];
// ----- Local connection due to Wire 176 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[17] = chanx_right_in[16];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[18] = chanx_right_in[17];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[19] = chanx_right_in[18];
// ----- Local connection due to Wire 180 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[21] = chanx_right_in[20];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[22] = chanx_right_in[21];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[23] = chanx_right_in[22];
// ----- Local connection due to Wire 184 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[25] = chanx_right_in[24];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[26] = chanx_right_in[25];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[27] = chanx_right_in[26];
// ----- Local connection due to Wire 188 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[29] = chanx_right_in[28];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[30] = chanx_right_in[29];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[31] = chanx_right_in[30];
// ----- Local connection due to Wire 192 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[33] = chanx_right_in[32];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[34] = chanx_right_in[33];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[35] = chanx_right_in[34];
// ----- Local connection due to Wire 196 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[37] = chanx_right_in[36];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[38] = chanx_right_in[37];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[39] = chanx_right_in[38];
// ----- Local connection due to Wire 200 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[41] = chanx_right_in[40];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[42] = chanx_right_in[41];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[43] = chanx_right_in[42];
// ----- Local connection due to Wire 204 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[45] = chanx_right_in[44];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[46] = chanx_right_in[45];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[47] = chanx_right_in[46];
// ----- Local connection due to Wire 208 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[49] = chanx_right_in[48];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[50] = chanx_right_in[49];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[51] = chanx_right_in[50];
// ----- Local connection due to Wire 212 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[53] = chanx_right_in[52];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[54] = chanx_right_in[53];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[55] = chanx_right_in[54];
// ----- Local connection due to Wire 216 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[57] = chanx_right_in[56];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[58] = chanx_right_in[57];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[59] = chanx_right_in[58];
// ----- Local connection due to Wire 220 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[61] = chanx_right_in[60];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[62] = chanx_right_in[61];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[63] = chanx_right_in[62];
// ----- Local connection due to Wire 224 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[65] = chanx_right_in[64];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[66] = chanx_right_in[65];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[67] = chanx_right_in[66];
// ----- Local connection due to Wire 228 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[69] = chanx_right_in[68];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[70] = chanx_right_in[69];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[71] = chanx_right_in[70];
// ----- Local connection due to Wire 232 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[73] = chanx_right_in[72];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[74] = chanx_right_in[73];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[75] = chanx_right_in[74];
// ----- Local connection due to Wire 236 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[77] = chanx_right_in[76];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[78] = chanx_right_in[77];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[79] = chanx_right_in[78];
// ----- Local connection due to Wire 240 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[81] = chanx_right_in[80];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[82] = chanx_right_in[81];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[83] = chanx_right_in[82];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[85] = chanx_right_in[84];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[86] = chanx_right_in[85];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[87] = chanx_right_in[86];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[89] = chanx_right_in[88];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[90] = chanx_right_in[89];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[91] = chanx_right_in[90];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[93] = chanx_right_in[92];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[94] = chanx_right_in[93];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[95] = chanx_right_in[94];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[97] = chanx_right_in[96];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[98] = chanx_right_in[97];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[99] = chanx_right_in[98];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[101] = chanx_right_in[100];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[102] = chanx_right_in[101];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 2 -----
	assign chanx_left_out[103] = chanx_right_in[102];
// ----- Local connection due to Wire 320 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 324 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 328 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 338 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 342 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 346 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 350 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 354 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 358 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 362 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 366 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 370 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 374 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 378 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 382 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 386 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 390 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 394 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 398 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 402 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 404 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 405 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 406 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 408 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 409 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 410 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 412 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 413 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 414 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 416 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 417 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 418 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 420 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 421 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 422 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 427 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[1] = chanx_left_in[0];
// ----- Local connection due to Wire 428 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[2] = chanx_left_in[1];
// ----- Local connection due to Wire 429 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[3] = chanx_left_in[2];
// ----- Local connection due to Wire 431 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[5] = chanx_left_in[4];
// ----- Local connection due to Wire 432 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[6] = chanx_left_in[5];
// ----- Local connection due to Wire 433 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[7] = chanx_left_in[6];
// ----- Local connection due to Wire 435 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[9] = chanx_left_in[8];
// ----- Local connection due to Wire 436 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[10] = chanx_left_in[9];
// ----- Local connection due to Wire 437 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[11] = chanx_left_in[10];
// ----- Local connection due to Wire 439 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[13] = chanx_left_in[12];
// ----- Local connection due to Wire 440 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[14] = chanx_left_in[13];
// ----- Local connection due to Wire 441 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[15] = chanx_left_in[14];
// ----- Local connection due to Wire 443 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[17] = chanx_left_in[16];
// ----- Local connection due to Wire 444 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[18] = chanx_left_in[17];
// ----- Local connection due to Wire 445 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[19] = chanx_left_in[18];
// ----- Local connection due to Wire 447 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[21] = chanx_left_in[20];
// ----- Local connection due to Wire 448 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[22] = chanx_left_in[21];
// ----- Local connection due to Wire 449 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[23] = chanx_left_in[22];
// ----- Local connection due to Wire 451 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[25] = chanx_left_in[24];
// ----- Local connection due to Wire 452 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[26] = chanx_left_in[25];
// ----- Local connection due to Wire 453 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[27] = chanx_left_in[26];
// ----- Local connection due to Wire 455 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[29] = chanx_left_in[28];
// ----- Local connection due to Wire 456 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[30] = chanx_left_in[29];
// ----- Local connection due to Wire 457 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[31] = chanx_left_in[30];
// ----- Local connection due to Wire 459 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[33] = chanx_left_in[32];
// ----- Local connection due to Wire 460 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[34] = chanx_left_in[33];
// ----- Local connection due to Wire 461 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[35] = chanx_left_in[34];
// ----- Local connection due to Wire 463 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[37] = chanx_left_in[36];
// ----- Local connection due to Wire 464 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[38] = chanx_left_in[37];
// ----- Local connection due to Wire 465 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[39] = chanx_left_in[38];
// ----- Local connection due to Wire 467 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[41] = chanx_left_in[40];
// ----- Local connection due to Wire 468 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[42] = chanx_left_in[41];
// ----- Local connection due to Wire 469 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[43] = chanx_left_in[42];
// ----- Local connection due to Wire 471 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[45] = chanx_left_in[44];
// ----- Local connection due to Wire 472 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[46] = chanx_left_in[45];
// ----- Local connection due to Wire 473 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[47] = chanx_left_in[46];
// ----- Local connection due to Wire 475 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[49] = chanx_left_in[48];
// ----- Local connection due to Wire 476 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[50] = chanx_left_in[49];
// ----- Local connection due to Wire 477 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[51] = chanx_left_in[50];
// ----- Local connection due to Wire 479 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[53] = chanx_left_in[52];
// ----- Local connection due to Wire 480 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[54] = chanx_left_in[53];
// ----- Local connection due to Wire 481 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[55] = chanx_left_in[54];
// ----- Local connection due to Wire 483 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[57] = chanx_left_in[56];
// ----- Local connection due to Wire 484 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[58] = chanx_left_in[57];
// ----- Local connection due to Wire 485 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[59] = chanx_left_in[58];
// ----- Local connection due to Wire 487 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[61] = chanx_left_in[60];
// ----- Local connection due to Wire 488 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[62] = chanx_left_in[61];
// ----- Local connection due to Wire 489 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[63] = chanx_left_in[62];
// ----- Local connection due to Wire 491 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[65] = chanx_left_in[64];
// ----- Local connection due to Wire 492 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[66] = chanx_left_in[65];
// ----- Local connection due to Wire 493 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[67] = chanx_left_in[66];
// ----- Local connection due to Wire 495 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[69] = chanx_left_in[68];
// ----- Local connection due to Wire 496 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[70] = chanx_left_in[69];
// ----- Local connection due to Wire 497 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[71] = chanx_left_in[70];
// ----- Local connection due to Wire 499 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[73] = chanx_left_in[72];
// ----- Local connection due to Wire 500 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[74] = chanx_left_in[73];
// ----- Local connection due to Wire 501 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[75] = chanx_left_in[74];
// ----- Local connection due to Wire 503 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[77] = chanx_left_in[76];
// ----- Local connection due to Wire 504 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[78] = chanx_left_in[77];
// ----- Local connection due to Wire 505 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[79] = chanx_left_in[78];
// ----- Local connection due to Wire 507 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[81] = chanx_left_in[80];
// ----- Local connection due to Wire 508 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[82] = chanx_left_in[81];
// ----- Local connection due to Wire 509 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[83] = chanx_left_in[82];
// ----- Local connection due to Wire 511 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[85] = chanx_left_in[84];
// ----- Local connection due to Wire 512 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[86] = chanx_left_in[85];
// ----- Local connection due to Wire 513 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[87] = chanx_left_in[86];
// ----- Local connection due to Wire 515 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[89] = chanx_left_in[88];
// ----- Local connection due to Wire 516 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[90] = chanx_left_in[89];
// ----- Local connection due to Wire 517 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[91] = chanx_left_in[90];
// ----- Local connection due to Wire 519 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[93] = chanx_left_in[92];
// ----- Local connection due to Wire 520 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[94] = chanx_left_in[93];
// ----- Local connection due to Wire 521 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[95] = chanx_left_in[94];
// ----- Local connection due to Wire 523 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[97] = chanx_left_in[96];
// ----- Local connection due to Wire 524 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[98] = chanx_left_in[97];
// ----- Local connection due to Wire 525 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[99] = chanx_left_in[98];
// ----- Local connection due to Wire 527 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[101] = chanx_left_in[100];
// ----- Local connection due to Wire 528 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[102] = chanx_left_in[101];
// ----- Local connection due to Wire 529 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chanx_right_out[103] = chanx_left_in[102];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size15 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[1], chanx_right_in[7], chanx_right_in[37], chanx_right_in[73], chanx_left_in[0], chanx_left_in[3], chanx_left_in[36], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size15_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_0_sram_inv[0:3]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size15 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[13], chanx_right_in[43], chanx_right_in[49], chanx_right_in[85], chanx_left_in[24], chanx_left_in[60], chanx_left_in[75], chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size15_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_1_sram_inv[0:3]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size15 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_34_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovalid_2_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_4_0_, chanx_right_in[25], chanx_right_in[61], chanx_right_in[79], chanx_right_in[97], chanx_left_in[12], chanx_left_in[39], chanx_left_in[48], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size15_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_2_sram_inv[0:3]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size15 mux_right_track_72 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[46], chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[21], chany_bottom_in[57], chany_bottom_in[67], chany_bottom_in[93]}),
		.sram(mux_tree_tapbuf_size15_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_3_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size15 mux_right_track_144 (
		.in({chany_top_in[22], chany_top_in[58], chany_top_in[71], chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[45], chany_bottom_in[81]}),
		.sram(mux_tree_tapbuf_size15_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size15_4_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size15_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_0_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_1_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_2_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_3_sram_inv[0:3]));

	mux_tree_tapbuf_size15_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size15_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size15_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size15_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13 mux_top_track_8 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[2], chanx_right_in[11], chanx_right_in[38], chanx_right_in[74], chanx_left_in[34], chanx_left_in[70], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size13 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_, chanx_right_in[4], chanx_right_in[15], chanx_right_in[40], chanx_right_in[76], chanx_left_in[33], chanx_left_in[69], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size13 mux_top_track_24 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_, chanx_right_in[5], chanx_right_in[19], chanx_right_in[41], chanx_right_in[77], chanx_left_in[32], chanx_left_in[68], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size13 mux_top_track_184 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[32], chanx_right_in[68], chanx_right_in[99], chanx_left_in[5], chanx_left_in[19], chanx_left_in[41], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size13 mux_top_track_192 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[33], chanx_right_in[69], chanx_right_in[103], chanx_left_in[4], chanx_left_in[15], chanx_left_in[40], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size13 mux_top_track_200 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_, chanx_right_in[34], chanx_right_in[70], chanx_right_in[104], chanx_left_in[2], chanx_left_in[11], chanx_left_in[38], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size13 mux_right_track_0 (
		.in({chany_top_in[34], chany_top_in[70], chany_top_in[104], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_1_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_2_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_3_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_0_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[33], chany_bottom_in[69], chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size13 mux_right_track_8 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[36], chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, chany_bottom_in[32], chany_bottom_in[68], chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size13 mux_right_track_200 (
		.in({chany_top_in[32], chany_top_in[68], chany_top_in[99], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_, chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[36], chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size13_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size14 mux_top_track_32 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, chanx_right_in[6], chanx_right_in[23], chanx_right_in[42], chanx_right_in[78], chanx_left_in[30], chanx_left_in[66], chanx_left_in[95], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size14 mux_top_track_40 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[44], chanx_right_in[80], chanx_left_in[29], chanx_left_in[65], chanx_left_in[91], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size14_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_1_sram_inv[0:3]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size14 mux_top_track_48 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[9], chanx_right_in[31], chanx_right_in[45], chanx_right_in[81], chanx_left_in[28], chanx_left_in[64], chanx_left_in[87], chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size14_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_2_sram_inv[0:3]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size14 mux_top_track_56 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_, chanx_right_in[10], chanx_right_in[35], chanx_right_in[46], chanx_right_in[82], chanx_left_in[26], chanx_left_in[62], chanx_left_in[83], chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size14_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_3_sram_inv[0:3]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size14 mux_top_track_64 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_, chanx_right_in[12], chanx_right_in[39], chanx_right_in[48], chanx_right_in[84], chanx_left_in[25], chanx_left_in[61], chanx_left_in[79], chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size14_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_4_sram_inv[0:3]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size14 mux_top_track_80 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[14], chanx_right_in[47], chanx_right_in[50], chanx_right_in[86], chanx_left_in[22], chanx_left_in[58], chanx_left_in[71], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size14_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_5_sram_inv[0:3]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size14 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_, chanx_right_in[16], chanx_right_in[51:52], chanx_right_in[88], chanx_left_in[21], chanx_left_in[57], chanx_left_in[67], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size14_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_6_sram_inv[0:3]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size14 mux_top_track_96 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_, chanx_right_in[17], chanx_right_in[53], chanx_right_in[55], chanx_right_in[89], chanx_left_in[20], chanx_left_in[56], chanx_left_in[63], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size14_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_7_sram_inv[0:3]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size14 mux_top_track_104 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, chanx_right_in[18], chanx_right_in[54], chanx_right_in[59], chanx_right_in[90], chanx_left_in[18], chanx_left_in[54], chanx_left_in[59], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size14_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_8_sram_inv[0:3]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size14 mux_top_track_112 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_18_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_19_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_20_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_1_0_, chanx_right_in[20], chanx_right_in[56], chanx_right_in[63], chanx_right_in[92], chanx_left_in[17], chanx_left_in[53], chanx_left_in[55], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size14_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_9_sram_inv[0:3]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size14 mux_top_track_120 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_22_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_23_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_24_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_ordy_3_0_, chanx_right_in[21], chanx_right_in[57], chanx_right_in[67], chanx_right_in[93], chanx_left_in[16], chanx_left_in[51:52], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size14_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_10_sram_inv[0:3]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size14 mux_top_track_128 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_26_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_27_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_28_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_0_0_, chanx_right_in[22], chanx_right_in[58], chanx_right_in[71], chanx_right_in[94], chanx_left_in[14], chanx_left_in[47], chanx_left_in[50], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size14_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_11_sram_inv[0:3]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size14 mux_top_track_136 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_, chanx_right_in[24], chanx_right_in[60], chanx_right_in[75], chanx_right_in[96], chanx_left_in[13], chanx_left_in[43], chanx_left_in[49], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size14_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_12_sram_inv[0:3]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size14 mux_top_track_152 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_2_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_3_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_4_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_ovch_1_0_, chanx_right_in[26], chanx_right_in[62], chanx_right_in[83], chanx_right_in[98], chanx_left_in[10], chanx_left_in[35], chanx_left_in[46], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size14_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_13_sram_inv[0:3]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size14 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_6_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_7_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_8_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_0_0_, chanx_right_in[28], chanx_right_in[64], chanx_right_in[87], chanx_right_in[100], chanx_left_in[9], chanx_left_in[31], chanx_left_in[45], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size14_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_14_sram_inv[0:3]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size14 mux_top_track_168 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_10_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_11_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_12_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_2_0_, chanx_right_in[29], chanx_right_in[65], chanx_right_in[91], chanx_right_in[101], chanx_left_in[8], chanx_left_in[27], chanx_left_in[44], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size14_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_15_sram_inv[0:3]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size14 mux_top_track_176 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_14_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_15_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_16_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_oack_4_0_, chanx_right_in[30], chanx_right_in[66], chanx_right_in[95], chanx_right_in[102], chanx_left_in[6], chanx_left_in[23], chanx_left_in[42], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size14_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_16_sram_inv[0:3]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size14 mux_top_track_208 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_odata_0_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_1_30_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_2_31_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_3_32_, top_right_grid_left_width_0_height_0_subtile_0__pin_odata_4_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_olck_2_0_, chanx_right_in[0], chanx_right_in[3], chanx_right_in[36], chanx_right_in[72], chanx_left_in[1], chanx_left_in[7], chanx_left_in[37], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_size14_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_17_sram_inv[0:3]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size14 mux_right_track_16 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[37], chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, chany_bottom_in[30], chany_bottom_in[66], chany_bottom_in[95], chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size14_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_18_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size14 mux_right_track_24 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[38], chany_top_in[74], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, chany_bottom_in[29], chany_bottom_in[65], chany_bottom_in[91], chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size14_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_19_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size14 mux_right_track_32 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[40], chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_, chany_bottom_in[28], chany_bottom_in[64], chany_bottom_in[87], chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size14_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_20_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size14 mux_right_track_40 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[41], chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[26], chany_bottom_in[62], chany_bottom_in[83], chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size14_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_21_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size14 mux_right_track_48 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[42], chany_top_in[78], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_, chany_bottom_in[25], chany_bottom_in[61], chany_bottom_in[79], chany_bottom_in[97]}),
		.sram(mux_tree_tapbuf_size14_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_22_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size14 mux_right_track_56 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[44], chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_, chany_bottom_in[24], chany_bottom_in[60], chany_bottom_in[75], chany_bottom_in[96]}),
		.sram(mux_tree_tapbuf_size14_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_23_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size14 mux_right_track_64 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[45], chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_, chany_bottom_in[22], chany_bottom_in[58], chany_bottom_in[71], chany_bottom_in[94]}),
		.sram(mux_tree_tapbuf_size14_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_24_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size14 mux_right_track_80 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[48], chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, chany_bottom_in[20], chany_bottom_in[56], chany_bottom_in[63], chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_size14_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_25_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size14 mux_right_track_88 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[49], chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, chany_bottom_in[18], chany_bottom_in[54], chany_bottom_in[59], chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size14_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_26_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size14 mux_right_track_96 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[50], chany_top_in[86], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, chany_bottom_in[17], chany_bottom_in[53], chany_bottom_in[55], chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_size14_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_27_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size14 mux_right_track_104 (
		.in({chany_top_in[16], chany_top_in[51:52], chany_top_in[88], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_, chany_bottom_in[16], chany_bottom_in[51:52], chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_size14_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_28_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size14 mux_right_track_112 (
		.in({chany_top_in[17], chany_top_in[53], chany_top_in[55], chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[50], chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_size14_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_29_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size14 mux_right_track_120 (
		.in({chany_top_in[18], chany_top_in[54], chany_top_in[59], chany_top_in[90], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_, chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[49], chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_size14_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_30_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size14 mux_right_track_128 (
		.in({chany_top_in[20], chany_top_in[56], chany_top_in[63], chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_29_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_30_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_31_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_1_1_, chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[48], chany_bottom_in[84]}),
		.sram(mux_tree_tapbuf_size14_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_31_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size14 mux_right_track_136 (
		.in({chany_top_in[21], chany_top_in[57], chany_top_in[67], chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_, chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[46], chany_bottom_in[82]}),
		.sram(mux_tree_tapbuf_size14_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_32_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size14 mux_right_track_152 (
		.in({chany_top_in[24], chany_top_in[60], chany_top_in[75], chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_5_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_6_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_7_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovch_4_0_, chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[44], chany_bottom_in[80]}),
		.sram(mux_tree_tapbuf_size14_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_33_sram_inv[0:3]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size14 mux_right_track_160 (
		.in({chany_top_in[25], chany_top_in[61], chany_top_in[79], chany_top_in[97], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_9_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_10_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_11_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_1_1_, chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[42], chany_bottom_in[78]}),
		.sram(mux_tree_tapbuf_size14_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_34_sram_inv[0:3]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size14 mux_right_track_168 (
		.in({chany_top_in[26], chany_top_in[62], chany_top_in[83], chany_top_in[98], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_13_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_14_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_15_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_oack_3_1_, chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[41], chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size14_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_35_sram_inv[0:3]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size14 mux_right_track_176 (
		.in({chany_top_in[28], chany_top_in[64], chany_top_in[87], chany_top_in[100], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_17_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_18_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_19_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_0_1_, chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[40], chany_bottom_in[76]}),
		.sram(mux_tree_tapbuf_size14_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_36_sram_inv[0:3]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size14 mux_right_track_184 (
		.in({chany_top_in[29], chany_top_in[65], chany_top_in[91], chany_top_in[101], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_21_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_22_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_23_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_2_1_, chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[38], chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_size14_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_37_sram_inv[0:3]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size14 mux_right_track_192 (
		.in({chany_top_in[30], chany_top_in[66], chany_top_in[95], chany_top_in[102], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_25_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_26_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_3_27_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ordy_4_1_, chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_size14_38_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_38_sram_inv[0:3]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size14_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_1_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_2_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_3_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_4_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_5_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_6_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_7_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_8_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_9_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_10_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_11_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_12_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_13_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_14_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_15_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_16_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_17_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_18_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_19_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_20_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_21_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_22_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_23_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_24_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_25_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_26_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_27_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_28_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_29_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_30_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_31_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_32_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size15_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_33_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_34_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_35_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_36_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_37_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_38_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_38_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_right_track_208 (
		.in({chany_top_in[33], chany_top_in[69], chany_top_in[103], right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_0_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_1_33_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_2_34_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_odata_4_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_ovalid_1_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_olck_3_1_, chany_bottom_in[34], chany_bottom_in[70], chany_bottom_in[104]}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size12_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size8 mux_bottom_track_1 (
		.in({chanx_right_in[33], chanx_right_in[69], chanx_right_in[103], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[1], chanx_left_in[7], chanx_left_in[37], chanx_left_in[73]}),
		.sram(mux_tree_tapbuf_size8_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_0_sram_inv[0:3]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size8 mux_bottom_track_9 (
		.in({chanx_right_in[32], chanx_right_in[68], chanx_right_in[99], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[2], chanx_left_in[11], chanx_left_in[38], chanx_left_in[74]}),
		.sram(mux_tree_tapbuf_size8_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_1_sram_inv[0:3]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size8 mux_bottom_track_17 (
		.in({chanx_right_in[30], chanx_right_in[66], chanx_right_in[95], chanx_right_in[102], chanx_left_in[4], chanx_left_in[15], chanx_left_in[40], chanx_left_in[76]}),
		.sram(mux_tree_tapbuf_size8_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_2_sram_inv[0:3]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size8 mux_bottom_track_25 (
		.in({chanx_right_in[29], chanx_right_in[65], chanx_right_in[91], chanx_right_in[101], chanx_left_in[5], chanx_left_in[19], chanx_left_in[41], chanx_left_in[77]}),
		.sram(mux_tree_tapbuf_size8_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_3_sram_inv[0:3]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size8 mux_bottom_track_33 (
		.in({chanx_right_in[28], chanx_right_in[64], chanx_right_in[87], chanx_right_in[100], chanx_left_in[6], chanx_left_in[23], chanx_left_in[42], chanx_left_in[78]}),
		.sram(mux_tree_tapbuf_size8_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_4_sram_inv[0:3]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size8 mux_bottom_track_41 (
		.in({chanx_right_in[26], chanx_right_in[62], chanx_right_in[83], chanx_right_in[98], chanx_left_in[8], chanx_left_in[27], chanx_left_in[44], chanx_left_in[80]}),
		.sram(mux_tree_tapbuf_size8_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_5_sram_inv[0:3]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size8 mux_bottom_track_49 (
		.in({chanx_right_in[25], chanx_right_in[61], chanx_right_in[79], chanx_right_in[97], chanx_left_in[9], chanx_left_in[31], chanx_left_in[45], chanx_left_in[81]}),
		.sram(mux_tree_tapbuf_size8_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_6_sram_inv[0:3]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size8 mux_bottom_track_57 (
		.in({chanx_right_in[24], chanx_right_in[60], chanx_right_in[75], chanx_right_in[96], chanx_left_in[10], chanx_left_in[35], chanx_left_in[46], chanx_left_in[82]}),
		.sram(mux_tree_tapbuf_size8_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_7_sram_inv[0:3]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size8 mux_bottom_track_65 (
		.in({chanx_right_in[22], chanx_right_in[58], chanx_right_in[71], chanx_right_in[94], chanx_left_in[12], chanx_left_in[39], chanx_left_in[48], chanx_left_in[84]}),
		.sram(mux_tree_tapbuf_size8_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_8_sram_inv[0:3]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size8 mux_bottom_track_89 (
		.in({chanx_right_in[18], chanx_right_in[54], chanx_right_in[59], chanx_right_in[90], chanx_left_in[16], chanx_left_in[51:52], chanx_left_in[88]}),
		.sram(mux_tree_tapbuf_size8_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_9_sram_inv[0:3]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size8 mux_bottom_track_97 (
		.in({chanx_right_in[17], chanx_right_in[53], chanx_right_in[55], chanx_right_in[89], chanx_left_in[17], chanx_left_in[53], chanx_left_in[55], chanx_left_in[89]}),
		.sram(mux_tree_tapbuf_size8_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_10_sram_inv[0:3]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size8 mux_bottom_track_105 (
		.in({chanx_right_in[16], chanx_right_in[51:52], chanx_right_in[88], chanx_left_in[18], chanx_left_in[54], chanx_left_in[59], chanx_left_in[90]}),
		.sram(mux_tree_tapbuf_size8_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_11_sram_inv[0:3]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size8 mux_bottom_track_113 (
		.in({chanx_right_in[14], chanx_right_in[47], chanx_right_in[50], chanx_right_in[86], chanx_left_in[20], chanx_left_in[56], chanx_left_in[63], chanx_left_in[92]}),
		.sram(mux_tree_tapbuf_size8_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_12_sram_inv[0:3]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size8 mux_bottom_track_121 (
		.in({chanx_right_in[13], chanx_right_in[43], chanx_right_in[49], chanx_right_in[85], chanx_left_in[21], chanx_left_in[57], chanx_left_in[67], chanx_left_in[93]}),
		.sram(mux_tree_tapbuf_size8_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_13_sram_inv[0:3]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size8 mux_bottom_track_129 (
		.in({chanx_right_in[12], chanx_right_in[39], chanx_right_in[48], chanx_right_in[84], chanx_left_in[22], chanx_left_in[58], chanx_left_in[71], chanx_left_in[94]}),
		.sram(mux_tree_tapbuf_size8_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_14_sram_inv[0:3]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size8 mux_bottom_track_137 (
		.in({chanx_right_in[10], chanx_right_in[35], chanx_right_in[46], chanx_right_in[82], chanx_left_in[24], chanx_left_in[60], chanx_left_in[75], chanx_left_in[96]}),
		.sram(mux_tree_tapbuf_size8_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_15_sram_inv[0:3]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size8 mux_bottom_track_161 (
		.in({chanx_right_in[6], chanx_right_in[23], chanx_right_in[42], chanx_right_in[78], chanx_left_in[28], chanx_left_in[64], chanx_left_in[87], chanx_left_in[100]}),
		.sram(mux_tree_tapbuf_size8_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_16_sram_inv[0:3]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size8 mux_bottom_track_169 (
		.in({chanx_right_in[5], chanx_right_in[19], chanx_right_in[41], chanx_right_in[77], chanx_left_in[29], chanx_left_in[65], chanx_left_in[91], chanx_left_in[101]}),
		.sram(mux_tree_tapbuf_size8_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_17_sram_inv[0:3]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size8 mux_bottom_track_177 (
		.in({chanx_right_in[4], chanx_right_in[15], chanx_right_in[40], chanx_right_in[76], chanx_left_in[30], chanx_left_in[66], chanx_left_in[95], chanx_left_in[102]}),
		.sram(mux_tree_tapbuf_size8_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_18_sram_inv[0:3]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size8 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], chany_top_in[36], chany_top_in[72], chany_bottom_in[34], chany_bottom_in[70], chany_bottom_in[104], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size8_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_19_sram_inv[0:3]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size8 mux_left_track_9 (
		.in({chany_top_in[34], chany_top_in[70], chany_top_in[104], chany_bottom_in[0], chany_bottom_in[3], chany_bottom_in[36], chany_bottom_in[72], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size8_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_20_sram_inv[0:3]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size8 mux_left_track_33 (
		.in({chany_top_in[30], chany_top_in[66], chany_top_in[95], chany_top_in[102], chany_bottom_in[4], chany_bottom_in[15], chany_bottom_in[40], chany_bottom_in[76]}),
		.sram(mux_tree_tapbuf_size8_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_21_sram_inv[0:3]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size8 mux_left_track_41 (
		.in({chany_top_in[29], chany_top_in[65], chany_top_in[91], chany_top_in[101], chany_bottom_in[5], chany_bottom_in[19], chany_bottom_in[41], chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size8_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_22_sram_inv[0:3]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size8 mux_left_track_49 (
		.in({chany_top_in[28], chany_top_in[64], chany_top_in[87], chany_top_in[100], chany_bottom_in[6], chany_bottom_in[23], chany_bottom_in[42], chany_bottom_in[78]}),
		.sram(mux_tree_tapbuf_size8_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_23_sram_inv[0:3]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size8 mux_left_track_57 (
		.in({chany_top_in[26], chany_top_in[62], chany_top_in[83], chany_top_in[98], chany_bottom_in[8], chany_bottom_in[27], chany_bottom_in[44], chany_bottom_in[80]}),
		.sram(mux_tree_tapbuf_size8_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_24_sram_inv[0:3]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size8 mux_left_track_65 (
		.in({chany_top_in[25], chany_top_in[61], chany_top_in[79], chany_top_in[97], chany_bottom_in[9], chany_bottom_in[31], chany_bottom_in[45], chany_bottom_in[81]}),
		.sram(mux_tree_tapbuf_size8_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_25_sram_inv[0:3]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size8 mux_left_track_89 (
		.in({chany_top_in[21], chany_top_in[57], chany_top_in[67], chany_top_in[93], chany_bottom_in[13], chany_bottom_in[43], chany_bottom_in[49], chany_bottom_in[85]}),
		.sram(mux_tree_tapbuf_size8_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_26_sram_inv[0:3]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size8 mux_left_track_97 (
		.in({chany_top_in[20], chany_top_in[56], chany_top_in[63], chany_top_in[92], chany_bottom_in[14], chany_bottom_in[47], chany_bottom_in[50], chany_bottom_in[86]}),
		.sram(mux_tree_tapbuf_size8_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_27_sram_inv[0:3]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size8 mux_left_track_105 (
		.in({chany_top_in[18], chany_top_in[54], chany_top_in[59], chany_top_in[90], chany_bottom_in[16], chany_bottom_in[51:52], chany_bottom_in[88]}),
		.sram(mux_tree_tapbuf_size8_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_28_sram_inv[0:3]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size8 mux_left_track_113 (
		.in({chany_top_in[17], chany_top_in[53], chany_top_in[55], chany_top_in[89], chany_bottom_in[17], chany_bottom_in[53], chany_bottom_in[55], chany_bottom_in[89]}),
		.sram(mux_tree_tapbuf_size8_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_29_sram_inv[0:3]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size8 mux_left_track_121 (
		.in({chany_top_in[16], chany_top_in[51:52], chany_top_in[88], chany_bottom_in[18], chany_bottom_in[54], chany_bottom_in[59], chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size8_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_30_sram_inv[0:3]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size8 mux_left_track_129 (
		.in({chany_top_in[14], chany_top_in[47], chany_top_in[50], chany_top_in[86], chany_bottom_in[20], chany_bottom_in[56], chany_bottom_in[63], chany_bottom_in[92]}),
		.sram(mux_tree_tapbuf_size8_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_31_sram_inv[0:3]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size8 mux_left_track_137 (
		.in({chany_top_in[13], chany_top_in[43], chany_top_in[49], chany_top_in[85], chany_bottom_in[21], chany_bottom_in[57], chany_bottom_in[67], chany_bottom_in[93]}),
		.sram(mux_tree_tapbuf_size8_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_32_sram_inv[0:3]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size8 mux_left_track_161 (
		.in({chany_top_in[9], chany_top_in[31], chany_top_in[45], chany_top_in[81], chany_bottom_in[25], chany_bottom_in[61], chany_bottom_in[79], chany_bottom_in[97]}),
		.sram(mux_tree_tapbuf_size8_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_33_sram_inv[0:3]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size8 mux_left_track_169 (
		.in({chany_top_in[8], chany_top_in[27], chany_top_in[44], chany_top_in[80], chany_bottom_in[26], chany_bottom_in[62], chany_bottom_in[83], chany_bottom_in[98]}),
		.sram(mux_tree_tapbuf_size8_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_34_sram_inv[0:3]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size8 mux_left_track_177 (
		.in({chany_top_in[6], chany_top_in[23], chany_top_in[42], chany_top_in[78], chany_bottom_in[28], chany_bottom_in[64], chany_bottom_in[87], chany_bottom_in[100]}),
		.sram(mux_tree_tapbuf_size8_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_35_sram_inv[0:3]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size8 mux_left_track_185 (
		.in({chany_top_in[5], chany_top_in[19], chany_top_in[41], chany_top_in[77], chany_bottom_in[29], chany_bottom_in[65], chany_bottom_in[91], chany_bottom_in[101]}),
		.sram(mux_tree_tapbuf_size8_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_36_sram_inv[0:3]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size8 mux_left_track_193 (
		.in({chany_top_in[4], chany_top_in[15], chany_top_in[40], chany_top_in[76], chany_bottom_in[30], chany_bottom_in[66], chany_bottom_in[95], chany_bottom_in[102]}),
		.sram(mux_tree_tapbuf_size8_37_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size8_37_sram_inv[0:3]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_0_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_1_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_2_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_3_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_4_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_5_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_6_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_7_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_8_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_9_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_10_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_11_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_12_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_13_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_14_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_15_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_16_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_17_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_18_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_19_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_20_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_21_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_22_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_23_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_24_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_25_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_26_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_27_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_28_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_29_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_30_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_31_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_32_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_33_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_34_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_35_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_36_sram_inv[0:3]));

	mux_tree_tapbuf_size8_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size8_37_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size8_37_sram_inv[0:3]));

	mux_tree_tapbuf_size9 mux_bottom_track_73 (
		.in({chanx_right_in[21], chanx_right_in[57], chanx_right_in[67], chanx_right_in[93], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[13], chanx_left_in[43], chanx_left_in[49], chanx_left_in[85]}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size9 mux_bottom_track_81 (
		.in({chanx_right_in[20], chanx_right_in[56], chanx_right_in[63], chanx_right_in[92], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[14], chanx_left_in[47], chanx_left_in[50], chanx_left_in[86]}),
		.sram(mux_tree_tapbuf_size9_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_1_sram_inv[0:3]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size9 mux_bottom_track_145 (
		.in({chanx_right_in[9], chanx_right_in[31], chanx_right_in[45], chanx_right_in[81], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_left_in[25], chanx_left_in[61], chanx_left_in[79], chanx_left_in[97]}),
		.sram(mux_tree_tapbuf_size9_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_2_sram_inv[0:3]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size9 mux_bottom_track_153 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[44], chanx_right_in[80], bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[26], chanx_left_in[62], chanx_left_in[83], chanx_left_in[98]}),
		.sram(mux_tree_tapbuf_size9_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_3_sram_inv[0:3]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size9 mux_left_track_73 (
		.in({chany_top_in[24], chany_top_in[60], chany_top_in[75], chany_top_in[96], chany_bottom_in[10], chany_bottom_in[35], chany_bottom_in[46], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_4_sram_inv[0:3]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size9 mux_left_track_81 (
		.in({chany_top_in[22], chany_top_in[58], chany_top_in[71], chany_top_in[94], chany_bottom_in[12], chany_bottom_in[39], chany_bottom_in[48], chany_bottom_in[84], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_5_sram_inv[0:3]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size9 mux_left_track_145 (
		.in({chany_top_in[12], chany_top_in[39], chany_top_in[48], chany_top_in[84], chany_bottom_in[22], chany_bottom_in[58], chany_bottom_in[71], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_}),
		.sram(mux_tree_tapbuf_size9_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_6_sram_inv[0:3]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size9 mux_left_track_153 (
		.in({chany_top_in[10], chany_top_in[35], chany_top_in[46], chany_top_in[82], chany_bottom_in[24], chany_bottom_in[60], chany_bottom_in[75], chany_bottom_in[96], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size9_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_7_sram_inv[0:3]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_1_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_2_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_3_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_4_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_5_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_6_sram_inv[0:3]));

	mux_tree_tapbuf_size9_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_7_sram_inv[0:3]));

	mux_tree_tapbuf_size7 mux_bottom_track_185 (
		.in({chanx_right_in[2], chanx_right_in[11], chanx_right_in[38], chanx_right_in[74], chanx_left_in[32], chanx_left_in[68], chanx_left_in[99]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size7 mux_bottom_track_193 (
		.in({chanx_right_in[1], chanx_right_in[7], chanx_right_in[37], chanx_right_in[73], chanx_left_in[33], chanx_left_in[69], chanx_left_in[103]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size7 mux_bottom_track_201 (
		.in({chanx_right_in[0], chanx_right_in[3], chanx_right_in[36], chanx_right_in[72], chanx_left_in[34], chanx_left_in[70], chanx_left_in[104]}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size7 mux_bottom_track_209 (
		.in({chanx_right_in[34], chanx_right_in[70], chanx_right_in[104], chanx_left_in[0], chanx_left_in[3], chanx_left_in[36], chanx_left_in[72]}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size7 mux_left_track_17 (
		.in({chany_top_in[33], chany_top_in[69], chany_top_in[103], chany_bottom_in[1], chany_bottom_in[7], chany_bottom_in[37], chany_bottom_in[73]}),
		.sram(mux_tree_tapbuf_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_4_sram_inv[0:2]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size7 mux_left_track_25 (
		.in({chany_top_in[32], chany_top_in[68], chany_top_in[99], chany_bottom_in[2], chany_bottom_in[11], chany_bottom_in[38], chany_bottom_in[74]}),
		.sram(mux_tree_tapbuf_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_5_sram_inv[0:2]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size7 mux_left_track_201 (
		.in({chany_top_in[2], chany_top_in[11], chany_top_in[38], chany_top_in[74], chany_bottom_in[32], chany_bottom_in[68], chany_bottom_in[99]}),
		.sram(mux_tree_tapbuf_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_6_sram_inv[0:2]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size7 mux_left_track_209 (
		.in({chany_top_in[1], chany_top_in[7], chany_top_in[37], chany_top_in[73], chany_bottom_in[33], chany_bottom_in[69], chany_bottom_in[103]}),
		.sram(mux_tree_tapbuf_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_7_sram_inv[0:2]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size8_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_7_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_5__5_ -----

//----- Default net type -----
`default_nettype wire



