//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: router_tb
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Jun 29 10:24:47 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

module router_tb_top_formal_verification (
input [0:0] clk,
input [0:0] reset,
input [0:0] channel_in_ip_67_,
input [0:0] channel_in_ip_66_,
input [0:0] channel_in_ip_65_,
input [0:0] channel_in_ip_64_,
input [0:0] channel_in_ip_63_,
input [0:0] channel_in_ip_62_,
input [0:0] channel_in_ip_61_,
input [0:0] channel_in_ip_60_,
input [0:0] channel_in_ip_59_,
input [0:0] channel_in_ip_58_,
input [0:0] channel_in_ip_57_,
input [0:0] channel_in_ip_56_,
input [0:0] channel_in_ip_55_,
input [0:0] channel_in_ip_54_,
input [0:0] channel_in_ip_53_,
input [0:0] channel_in_ip_52_,
input [0:0] channel_in_ip_51_,
input [0:0] channel_in_ip_50_,
input [0:0] channel_in_ip_49_,
input [0:0] channel_in_ip_48_,
input [0:0] channel_in_ip_47_,
input [0:0] channel_in_ip_46_,
input [0:0] channel_in_ip_45_,
input [0:0] channel_in_ip_44_,
input [0:0] channel_in_ip_43_,
input [0:0] channel_in_ip_42_,
input [0:0] channel_in_ip_41_,
input [0:0] channel_in_ip_40_,
input [0:0] channel_in_ip_39_,
input [0:0] channel_in_ip_38_,
input [0:0] channel_in_ip_37_,
input [0:0] channel_in_ip_36_,
input [0:0] channel_in_ip_35_,
input [0:0] channel_in_ip_34_,
input [0:0] channel_in_ip_33_,
input [0:0] channel_in_ip_32_,
input [0:0] channel_in_ip_31_,
input [0:0] channel_in_ip_30_,
input [0:0] channel_in_ip_29_,
input [0:0] channel_in_ip_28_,
input [0:0] channel_in_ip_27_,
input [0:0] channel_in_ip_26_,
input [0:0] channel_in_ip_25_,
input [0:0] channel_in_ip_24_,
input [0:0] channel_in_ip_23_,
input [0:0] channel_in_ip_22_,
input [0:0] channel_in_ip_21_,
input [0:0] channel_in_ip_20_,
input [0:0] channel_in_ip_19_,
input [0:0] channel_in_ip_18_,
input [0:0] channel_in_ip_17_,
input [0:0] channel_in_ip_16_,
input [0:0] channel_in_ip_15_,
input [0:0] channel_in_ip_14_,
input [0:0] channel_in_ip_13_,
input [0:0] channel_in_ip_12_,
input [0:0] channel_in_ip_11_,
input [0:0] channel_in_ip_10_,
input [0:0] channel_in_ip_9_,
input [0:0] channel_in_ip_8_,
input [0:0] channel_in_ip_7_,
input [0:0] channel_in_ip_6_,
input [0:0] channel_in_ip_5_,
input [0:0] channel_in_ip_4_,
input [0:0] channel_in_ip_3_,
input [0:0] channel_in_ip_2_,
input [0:0] channel_in_ip_1_,
input [0:0] channel_in_ip_0_,
output [0:0] channel_out_op_67_,
output [0:0] channel_out_op_66_,
output [0:0] channel_out_op_65_,
output [0:0] channel_out_op_64_,
output [0:0] channel_out_op_63_,
output [0:0] channel_out_op_62_,
output [0:0] channel_out_op_61_,
output [0:0] channel_out_op_60_,
output [0:0] channel_out_op_59_,
output [0:0] channel_out_op_58_,
output [0:0] channel_out_op_57_,
output [0:0] channel_out_op_56_,
output [0:0] channel_out_op_55_,
output [0:0] channel_out_op_54_,
output [0:0] channel_out_op_53_,
output [0:0] channel_out_op_52_,
output [0:0] channel_out_op_51_,
output [0:0] channel_out_op_50_,
output [0:0] channel_out_op_49_,
output [0:0] channel_out_op_48_,
output [0:0] channel_out_op_47_,
output [0:0] channel_out_op_46_,
output [0:0] channel_out_op_45_,
output [0:0] channel_out_op_44_,
output [0:0] channel_out_op_43_,
output [0:0] channel_out_op_42_,
output [0:0] channel_out_op_41_,
output [0:0] channel_out_op_40_,
output [0:0] channel_out_op_39_,
output [0:0] channel_out_op_38_,
output [0:0] channel_out_op_37_,
output [0:0] channel_out_op_36_,
output [0:0] channel_out_op_35_,
output [0:0] channel_out_op_34_,
output [0:0] channel_out_op_33_,
output [0:0] channel_out_op_32_,
output [0:0] channel_out_op_31_,
output [0:0] channel_out_op_30_,
output [0:0] channel_out_op_29_,
output [0:0] channel_out_op_28_,
output [0:0] channel_out_op_27_,
output [0:0] channel_out_op_26_,
output [0:0] channel_out_op_25_,
output [0:0] channel_out_op_24_,
output [0:0] channel_out_op_23_,
output [0:0] channel_out_op_22_,
output [0:0] channel_out_op_21_,
output [0:0] channel_out_op_20_,
output [0:0] channel_out_op_19_,
output [0:0] channel_out_op_18_,
output [0:0] channel_out_op_17_,
output [0:0] channel_out_op_16_,
output [0:0] channel_out_op_15_,
output [0:0] channel_out_op_14_,
output [0:0] channel_out_op_13_,
output [0:0] channel_out_op_12_,
output [0:0] channel_out_op_11_,
output [0:0] channel_out_op_10_,
output [0:0] channel_out_op_9_,
output [0:0] channel_out_op_8_,
output [0:0] channel_out_op_7_,
output [0:0] channel_out_op_6_,
output [0:0] channel_out_op_5_,
output [0:0] channel_out_op_4_,
output [0:0] channel_out_op_3_,
output [0:0] channel_out_op_2_,
output [0:0] channel_out_op_1_,
output [0:0] channel_out_op_0_,
output [0:0] rtr_error);

// ----- Local wires for FPGA fabric -----
wire [0:159] gfpga_pad_GPIO_PAD_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] prog_clk_fm;
wire [0:0] set_fm;
wire [0:0] reset_fm;
wire [0:0] clk_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		prog_clk_fm[0],
		set_fm[0],
		reset_fm[0],
		clk_fm[0],
		gfpga_pad_GPIO_PAD_fm[0:159],
		ccff_head_fm[0],
		ccff_tail_fm[0]);

// ----- Begin Connect Global ports of FPGA top module -----
	assign set_fm[0] = 1'b0;
	assign reset_fm[0] = 1'b0;
	assign clk_fm[0] = clk[0];
	assign prog_clk_fm[0] = 1'b0;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input clk is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[12] -----
	assign gfpga_pad_GPIO_PAD_fm[12] = clk[0];

// ----- Blif Benchmark input reset is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[88] -----
	assign gfpga_pad_GPIO_PAD_fm[88] = reset[0];

// ----- Blif Benchmark input channel_in_ip_67_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[119] -----
	assign gfpga_pad_GPIO_PAD_fm[119] = channel_in_ip_67_[0];

// ----- Blif Benchmark input channel_in_ip_66_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[113] -----
	assign gfpga_pad_GPIO_PAD_fm[113] = channel_in_ip_66_[0];

// ----- Blif Benchmark input channel_in_ip_65_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[130] -----
	assign gfpga_pad_GPIO_PAD_fm[130] = channel_in_ip_65_[0];

// ----- Blif Benchmark input channel_in_ip_64_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[111] -----
	assign gfpga_pad_GPIO_PAD_fm[111] = channel_in_ip_64_[0];

// ----- Blif Benchmark input channel_in_ip_63_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[139] -----
	assign gfpga_pad_GPIO_PAD_fm[139] = channel_in_ip_63_[0];

// ----- Blif Benchmark input channel_in_ip_62_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[148] -----
	assign gfpga_pad_GPIO_PAD_fm[148] = channel_in_ip_62_[0];

// ----- Blif Benchmark input channel_in_ip_61_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[116] -----
	assign gfpga_pad_GPIO_PAD_fm[116] = channel_in_ip_61_[0];

// ----- Blif Benchmark input channel_in_ip_60_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[117] -----
	assign gfpga_pad_GPIO_PAD_fm[117] = channel_in_ip_60_[0];

// ----- Blif Benchmark input channel_in_ip_59_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[136] -----
	assign gfpga_pad_GPIO_PAD_fm[136] = channel_in_ip_59_[0];

// ----- Blif Benchmark input channel_in_ip_58_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[141] -----
	assign gfpga_pad_GPIO_PAD_fm[141] = channel_in_ip_58_[0];

// ----- Blif Benchmark input channel_in_ip_57_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[101] -----
	assign gfpga_pad_GPIO_PAD_fm[101] = channel_in_ip_57_[0];

// ----- Blif Benchmark input channel_in_ip_56_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[7] -----
	assign gfpga_pad_GPIO_PAD_fm[7] = channel_in_ip_56_[0];

// ----- Blif Benchmark input channel_in_ip_55_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[135] -----
	assign gfpga_pad_GPIO_PAD_fm[135] = channel_in_ip_55_[0];

// ----- Blif Benchmark input channel_in_ip_54_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[147] -----
	assign gfpga_pad_GPIO_PAD_fm[147] = channel_in_ip_54_[0];

// ----- Blif Benchmark input channel_in_ip_53_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[153] -----
	assign gfpga_pad_GPIO_PAD_fm[153] = channel_in_ip_53_[0];

// ----- Blif Benchmark input channel_in_ip_52_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[1] -----
	assign gfpga_pad_GPIO_PAD_fm[1] = channel_in_ip_52_[0];

// ----- Blif Benchmark input channel_in_ip_51_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[2] -----
	assign gfpga_pad_GPIO_PAD_fm[2] = channel_in_ip_51_[0];

// ----- Blif Benchmark input channel_in_ip_50_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[152] -----
	assign gfpga_pad_GPIO_PAD_fm[152] = channel_in_ip_50_[0];

// ----- Blif Benchmark input channel_in_ip_49_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[134] -----
	assign gfpga_pad_GPIO_PAD_fm[134] = channel_in_ip_49_[0];

// ----- Blif Benchmark input channel_in_ip_48_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[127] -----
	assign gfpga_pad_GPIO_PAD_fm[127] = channel_in_ip_48_[0];

// ----- Blif Benchmark input channel_in_ip_47_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[159] -----
	assign gfpga_pad_GPIO_PAD_fm[159] = channel_in_ip_47_[0];

// ----- Blif Benchmark input channel_in_ip_46_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[126] -----
	assign gfpga_pad_GPIO_PAD_fm[126] = channel_in_ip_46_[0];

// ----- Blif Benchmark input channel_in_ip_45_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[142] -----
	assign gfpga_pad_GPIO_PAD_fm[142] = channel_in_ip_45_[0];

// ----- Blif Benchmark input channel_in_ip_44_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[4] -----
	assign gfpga_pad_GPIO_PAD_fm[4] = channel_in_ip_44_[0];

// ----- Blif Benchmark input channel_in_ip_43_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[157] -----
	assign gfpga_pad_GPIO_PAD_fm[157] = channel_in_ip_43_[0];

// ----- Blif Benchmark input channel_in_ip_42_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[132] -----
	assign gfpga_pad_GPIO_PAD_fm[132] = channel_in_ip_42_[0];

// ----- Blif Benchmark input channel_in_ip_41_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[121] -----
	assign gfpga_pad_GPIO_PAD_fm[121] = channel_in_ip_41_[0];

// ----- Blif Benchmark input channel_in_ip_40_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[114] -----
	assign gfpga_pad_GPIO_PAD_fm[114] = channel_in_ip_40_[0];

// ----- Blif Benchmark input channel_in_ip_39_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[104] -----
	assign gfpga_pad_GPIO_PAD_fm[104] = channel_in_ip_39_[0];

// ----- Blif Benchmark input channel_in_ip_38_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[5] -----
	assign gfpga_pad_GPIO_PAD_fm[5] = channel_in_ip_38_[0];

// ----- Blif Benchmark input channel_in_ip_37_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[156] -----
	assign gfpga_pad_GPIO_PAD_fm[156] = channel_in_ip_37_[0];

// ----- Blif Benchmark input channel_in_ip_36_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[6] -----
	assign gfpga_pad_GPIO_PAD_fm[6] = channel_in_ip_36_[0];

// ----- Blif Benchmark input channel_in_ip_35_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[129] -----
	assign gfpga_pad_GPIO_PAD_fm[129] = channel_in_ip_35_[0];

// ----- Blif Benchmark input channel_in_ip_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[151] -----
	assign gfpga_pad_GPIO_PAD_fm[151] = channel_in_ip_34_[0];

// ----- Blif Benchmark input channel_in_ip_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[144] -----
	assign gfpga_pad_GPIO_PAD_fm[144] = channel_in_ip_33_[0];

// ----- Blif Benchmark input channel_in_ip_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[120] -----
	assign gfpga_pad_GPIO_PAD_fm[120] = channel_in_ip_32_[0];

// ----- Blif Benchmark input channel_in_ip_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[109] -----
	assign gfpga_pad_GPIO_PAD_fm[109] = channel_in_ip_31_[0];

// ----- Blif Benchmark input channel_in_ip_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[110] -----
	assign gfpga_pad_GPIO_PAD_fm[110] = channel_in_ip_30_[0];

// ----- Blif Benchmark input channel_in_ip_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[149] -----
	assign gfpga_pad_GPIO_PAD_fm[149] = channel_in_ip_29_[0];

// ----- Blif Benchmark input channel_in_ip_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[146] -----
	assign gfpga_pad_GPIO_PAD_fm[146] = channel_in_ip_28_[0];

// ----- Blif Benchmark input channel_in_ip_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[97] -----
	assign gfpga_pad_GPIO_PAD_fm[97] = channel_in_ip_27_[0];

// ----- Blif Benchmark input channel_in_ip_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[106] -----
	assign gfpga_pad_GPIO_PAD_fm[106] = channel_in_ip_26_[0];

// ----- Blif Benchmark input channel_in_ip_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[158] -----
	assign gfpga_pad_GPIO_PAD_fm[158] = channel_in_ip_25_[0];

// ----- Blif Benchmark input channel_in_ip_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[112] -----
	assign gfpga_pad_GPIO_PAD_fm[112] = channel_in_ip_24_[0];

// ----- Blif Benchmark input channel_in_ip_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[115] -----
	assign gfpga_pad_GPIO_PAD_fm[115] = channel_in_ip_23_[0];

// ----- Blif Benchmark input channel_in_ip_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[145] -----
	assign gfpga_pad_GPIO_PAD_fm[145] = channel_in_ip_22_[0];

// ----- Blif Benchmark input channel_in_ip_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[138] -----
	assign gfpga_pad_GPIO_PAD_fm[138] = channel_in_ip_21_[0];

// ----- Blif Benchmark input channel_in_ip_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[143] -----
	assign gfpga_pad_GPIO_PAD_fm[143] = channel_in_ip_20_[0];

// ----- Blif Benchmark input channel_in_ip_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[3] -----
	assign gfpga_pad_GPIO_PAD_fm[3] = channel_in_ip_19_[0];

// ----- Blif Benchmark input channel_in_ip_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[150] -----
	assign gfpga_pad_GPIO_PAD_fm[150] = channel_in_ip_18_[0];

// ----- Blif Benchmark input channel_in_ip_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[128] -----
	assign gfpga_pad_GPIO_PAD_fm[128] = channel_in_ip_17_[0];

// ----- Blif Benchmark input channel_in_ip_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[118] -----
	assign gfpga_pad_GPIO_PAD_fm[118] = channel_in_ip_16_[0];

// ----- Blif Benchmark input channel_in_ip_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[131] -----
	assign gfpga_pad_GPIO_PAD_fm[131] = channel_in_ip_15_[0];

// ----- Blif Benchmark input channel_in_ip_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[137] -----
	assign gfpga_pad_GPIO_PAD_fm[137] = channel_in_ip_14_[0];

// ----- Blif Benchmark input channel_in_ip_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[11] -----
	assign gfpga_pad_GPIO_PAD_fm[11] = channel_in_ip_13_[0];

// ----- Blif Benchmark input channel_in_ip_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[124] -----
	assign gfpga_pad_GPIO_PAD_fm[124] = channel_in_ip_12_[0];

// ----- Blif Benchmark input channel_in_ip_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[107] -----
	assign gfpga_pad_GPIO_PAD_fm[107] = channel_in_ip_11_[0];

// ----- Blif Benchmark input channel_in_ip_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[108] -----
	assign gfpga_pad_GPIO_PAD_fm[108] = channel_in_ip_10_[0];

// ----- Blif Benchmark input channel_in_ip_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[123] -----
	assign gfpga_pad_GPIO_PAD_fm[123] = channel_in_ip_9_[0];

// ----- Blif Benchmark input channel_in_ip_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[122] -----
	assign gfpga_pad_GPIO_PAD_fm[122] = channel_in_ip_8_[0];

// ----- Blif Benchmark input channel_in_ip_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[105] -----
	assign gfpga_pad_GPIO_PAD_fm[105] = channel_in_ip_7_[0];

// ----- Blif Benchmark input channel_in_ip_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[125] -----
	assign gfpga_pad_GPIO_PAD_fm[125] = channel_in_ip_6_[0];

// ----- Blif Benchmark input channel_in_ip_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[13] -----
	assign gfpga_pad_GPIO_PAD_fm[13] = channel_in_ip_5_[0];

// ----- Blif Benchmark input channel_in_ip_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[8] -----
	assign gfpga_pad_GPIO_PAD_fm[8] = channel_in_ip_4_[0];

// ----- Blif Benchmark input channel_in_ip_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[140] -----
	assign gfpga_pad_GPIO_PAD_fm[140] = channel_in_ip_3_[0];

// ----- Blif Benchmark input channel_in_ip_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[154] -----
	assign gfpga_pad_GPIO_PAD_fm[154] = channel_in_ip_2_[0];

// ----- Blif Benchmark input channel_in_ip_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[14] -----
	assign gfpga_pad_GPIO_PAD_fm[14] = channel_in_ip_1_[0];

// ----- Blif Benchmark input channel_in_ip_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[133] -----
	assign gfpga_pad_GPIO_PAD_fm[133] = channel_in_ip_0_[0];

// ----- Blif Benchmark output channel_out_op_67_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[38] -----
	assign channel_out_op_67_[0] = gfpga_pad_GPIO_PAD_fm[38];

// ----- Blif Benchmark output channel_out_op_66_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[55] -----
	assign channel_out_op_66_[0] = gfpga_pad_GPIO_PAD_fm[55];

// ----- Blif Benchmark output channel_out_op_65_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[44] -----
	assign channel_out_op_65_[0] = gfpga_pad_GPIO_PAD_fm[44];

// ----- Blif Benchmark output channel_out_op_64_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[52] -----
	assign channel_out_op_64_[0] = gfpga_pad_GPIO_PAD_fm[52];

// ----- Blif Benchmark output channel_out_op_63_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[60] -----
	assign channel_out_op_63_[0] = gfpga_pad_GPIO_PAD_fm[60];

// ----- Blif Benchmark output channel_out_op_62_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[66] -----
	assign channel_out_op_62_[0] = gfpga_pad_GPIO_PAD_fm[66];

// ----- Blif Benchmark output channel_out_op_61_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[56] -----
	assign channel_out_op_61_[0] = gfpga_pad_GPIO_PAD_fm[56];

// ----- Blif Benchmark output channel_out_op_60_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[62] -----
	assign channel_out_op_60_[0] = gfpga_pad_GPIO_PAD_fm[62];

// ----- Blif Benchmark output channel_out_op_59_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[50] -----
	assign channel_out_op_59_[0] = gfpga_pad_GPIO_PAD_fm[50];

// ----- Blif Benchmark output channel_out_op_58_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[63] -----
	assign channel_out_op_58_[0] = gfpga_pad_GPIO_PAD_fm[63];

// ----- Blif Benchmark output channel_out_op_57_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[37] -----
	assign channel_out_op_57_[0] = gfpga_pad_GPIO_PAD_fm[37];

// ----- Blif Benchmark output channel_out_op_56_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[42] -----
	assign channel_out_op_56_[0] = gfpga_pad_GPIO_PAD_fm[42];

// ----- Blif Benchmark output channel_out_op_55_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[95] -----
	assign channel_out_op_55_[0] = gfpga_pad_GPIO_PAD_fm[95];

// ----- Blif Benchmark output channel_out_op_54_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[45] -----
	assign channel_out_op_54_[0] = gfpga_pad_GPIO_PAD_fm[45];

// ----- Blif Benchmark output channel_out_op_53_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[91] -----
	assign channel_out_op_53_[0] = gfpga_pad_GPIO_PAD_fm[91];

// ----- Blif Benchmark output channel_out_op_52_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[65] -----
	assign channel_out_op_52_[0] = gfpga_pad_GPIO_PAD_fm[65];

// ----- Blif Benchmark output channel_out_op_51_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[36] -----
	assign channel_out_op_51_[0] = gfpga_pad_GPIO_PAD_fm[36];

// ----- Blif Benchmark output channel_out_op_50_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[89] -----
	assign channel_out_op_50_[0] = gfpga_pad_GPIO_PAD_fm[89];

// ----- Blif Benchmark output channel_out_op_49_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[99] -----
	assign channel_out_op_49_[0] = gfpga_pad_GPIO_PAD_fm[99];

// ----- Blif Benchmark output channel_out_op_48_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[86] -----
	assign channel_out_op_48_[0] = gfpga_pad_GPIO_PAD_fm[86];

// ----- Blif Benchmark output channel_out_op_47_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[59] -----
	assign channel_out_op_47_[0] = gfpga_pad_GPIO_PAD_fm[59];

// ----- Blif Benchmark output channel_out_op_46_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[64] -----
	assign channel_out_op_46_[0] = gfpga_pad_GPIO_PAD_fm[64];

// ----- Blif Benchmark output channel_out_op_45_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[84] -----
	assign channel_out_op_45_[0] = gfpga_pad_GPIO_PAD_fm[84];

// ----- Blif Benchmark output channel_out_op_44_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[35] -----
	assign channel_out_op_44_[0] = gfpga_pad_GPIO_PAD_fm[35];

// ----- Blif Benchmark output channel_out_op_43_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[78] -----
	assign channel_out_op_43_[0] = gfpga_pad_GPIO_PAD_fm[78];

// ----- Blif Benchmark output channel_out_op_42_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[58] -----
	assign channel_out_op_42_[0] = gfpga_pad_GPIO_PAD_fm[58];

// ----- Blif Benchmark output channel_out_op_41_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[77] -----
	assign channel_out_op_41_[0] = gfpga_pad_GPIO_PAD_fm[77];

// ----- Blif Benchmark output channel_out_op_40_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[53] -----
	assign channel_out_op_40_[0] = gfpga_pad_GPIO_PAD_fm[53];

// ----- Blif Benchmark output channel_out_op_39_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[73] -----
	assign channel_out_op_39_[0] = gfpga_pad_GPIO_PAD_fm[73];

// ----- Blif Benchmark output channel_out_op_38_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[74] -----
	assign channel_out_op_38_[0] = gfpga_pad_GPIO_PAD_fm[74];

// ----- Blif Benchmark output channel_out_op_37_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[103] -----
	assign channel_out_op_37_[0] = gfpga_pad_GPIO_PAD_fm[103];

// ----- Blif Benchmark output channel_out_op_36_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[43] -----
	assign channel_out_op_36_[0] = gfpga_pad_GPIO_PAD_fm[43];

// ----- Blif Benchmark output channel_out_op_35_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[34] -----
	assign channel_out_op_35_[0] = gfpga_pad_GPIO_PAD_fm[34];

// ----- Blif Benchmark output channel_out_op_34_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[81] -----
	assign channel_out_op_34_[0] = gfpga_pad_GPIO_PAD_fm[81];

// ----- Blif Benchmark output channel_out_op_33_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[80] -----
	assign channel_out_op_33_[0] = gfpga_pad_GPIO_PAD_fm[80];

// ----- Blif Benchmark output channel_out_op_32_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[47] -----
	assign channel_out_op_32_[0] = gfpga_pad_GPIO_PAD_fm[47];

// ----- Blif Benchmark output channel_out_op_31_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[100] -----
	assign channel_out_op_31_[0] = gfpga_pad_GPIO_PAD_fm[100];

// ----- Blif Benchmark output channel_out_op_30_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[94] -----
	assign channel_out_op_30_[0] = gfpga_pad_GPIO_PAD_fm[94];

// ----- Blif Benchmark output channel_out_op_29_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[48] -----
	assign channel_out_op_29_[0] = gfpga_pad_GPIO_PAD_fm[48];

// ----- Blif Benchmark output channel_out_op_28_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[70] -----
	assign channel_out_op_28_[0] = gfpga_pad_GPIO_PAD_fm[70];

// ----- Blif Benchmark output channel_out_op_27_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[51] -----
	assign channel_out_op_27_[0] = gfpga_pad_GPIO_PAD_fm[51];

// ----- Blif Benchmark output channel_out_op_26_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[76] -----
	assign channel_out_op_26_[0] = gfpga_pad_GPIO_PAD_fm[76];

// ----- Blif Benchmark output channel_out_op_25_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[96] -----
	assign channel_out_op_25_[0] = gfpga_pad_GPIO_PAD_fm[96];

// ----- Blif Benchmark output channel_out_op_24_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[87] -----
	assign channel_out_op_24_[0] = gfpga_pad_GPIO_PAD_fm[87];

// ----- Blif Benchmark output channel_out_op_23_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[40] -----
	assign channel_out_op_23_[0] = gfpga_pad_GPIO_PAD_fm[40];

// ----- Blif Benchmark output channel_out_op_22_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[39] -----
	assign channel_out_op_22_[0] = gfpga_pad_GPIO_PAD_fm[39];

// ----- Blif Benchmark output channel_out_op_21_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[83] -----
	assign channel_out_op_21_[0] = gfpga_pad_GPIO_PAD_fm[83];

// ----- Blif Benchmark output channel_out_op_20_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[33] -----
	assign channel_out_op_20_[0] = gfpga_pad_GPIO_PAD_fm[33];

// ----- Blif Benchmark output channel_out_op_19_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[69] -----
	assign channel_out_op_19_[0] = gfpga_pad_GPIO_PAD_fm[69];

// ----- Blif Benchmark output channel_out_op_18_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[82] -----
	assign channel_out_op_18_[0] = gfpga_pad_GPIO_PAD_fm[82];

// ----- Blif Benchmark output channel_out_op_17_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[57] -----
	assign channel_out_op_17_[0] = gfpga_pad_GPIO_PAD_fm[57];

// ----- Blif Benchmark output channel_out_op_16_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[54] -----
	assign channel_out_op_16_[0] = gfpga_pad_GPIO_PAD_fm[54];

// ----- Blif Benchmark output channel_out_op_15_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[32] -----
	assign channel_out_op_15_[0] = gfpga_pad_GPIO_PAD_fm[32];

// ----- Blif Benchmark output channel_out_op_14_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[61] -----
	assign channel_out_op_14_[0] = gfpga_pad_GPIO_PAD_fm[61];

// ----- Blif Benchmark output channel_out_op_13_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[72] -----
	assign channel_out_op_13_[0] = gfpga_pad_GPIO_PAD_fm[72];

// ----- Blif Benchmark output channel_out_op_12_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[49] -----
	assign channel_out_op_12_[0] = gfpga_pad_GPIO_PAD_fm[49];

// ----- Blif Benchmark output channel_out_op_11_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[67] -----
	assign channel_out_op_11_[0] = gfpga_pad_GPIO_PAD_fm[67];

// ----- Blif Benchmark output channel_out_op_10_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[75] -----
	assign channel_out_op_10_[0] = gfpga_pad_GPIO_PAD_fm[75];

// ----- Blif Benchmark output channel_out_op_9_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[41] -----
	assign channel_out_op_9_[0] = gfpga_pad_GPIO_PAD_fm[41];

// ----- Blif Benchmark output channel_out_op_8_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[102] -----
	assign channel_out_op_8_[0] = gfpga_pad_GPIO_PAD_fm[102];

// ----- Blif Benchmark output channel_out_op_7_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[85] -----
	assign channel_out_op_7_[0] = gfpga_pad_GPIO_PAD_fm[85];

// ----- Blif Benchmark output channel_out_op_6_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[46] -----
	assign channel_out_op_6_[0] = gfpga_pad_GPIO_PAD_fm[46];

// ----- Blif Benchmark output channel_out_op_5_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[92] -----
	assign channel_out_op_5_[0] = gfpga_pad_GPIO_PAD_fm[92];

// ----- Blif Benchmark output channel_out_op_4_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[68] -----
	assign channel_out_op_4_[0] = gfpga_pad_GPIO_PAD_fm[68];

// ----- Blif Benchmark output channel_out_op_3_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[90] -----
	assign channel_out_op_3_[0] = gfpga_pad_GPIO_PAD_fm[90];

// ----- Blif Benchmark output channel_out_op_2_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[79] -----
	assign channel_out_op_2_[0] = gfpga_pad_GPIO_PAD_fm[79];

// ----- Blif Benchmark output channel_out_op_1_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[71] -----
	assign channel_out_op_1_[0] = gfpga_pad_GPIO_PAD_fm[71];

// ----- Blif Benchmark output channel_out_op_0_ is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[98] -----
	assign channel_out_op_0_[0] = gfpga_pad_GPIO_PAD_fm[98];

// ----- Blif Benchmark output rtr_error is mapped to FPGA IOPAD gfpga_pad_GPIO_PAD_fm[93] -----
	assign rtr_error[0] = gfpga_pad_GPIO_PAD_fm[93];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_GPIO_PAD_fm[0] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[9] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[10] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[15] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[16] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[17] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[18] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[19] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[20] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[21] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[22] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[23] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[24] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[25] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[26] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[27] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[28] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[29] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[30] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[31] = 1'b0;
	assign gfpga_pad_GPIO_PAD_fm[155] = 1'b0;

// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = 16'b1111111111001100;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = 16'b0000000000110011;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_out[0:15] = {16{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_mode_default__lut4_0.lut4_DFF_mem.mem_outb[0:15] = {16{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_n1_lut4__ble4_0.mem_ble4_out_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_0_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_1_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_2_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.mem_fle_3_in_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_1__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_2__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_3__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_4__7_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_5__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_4__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_3__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_2__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_1__0_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__1_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__2_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__3_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__4_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__5_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_0__6_.logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_DFF_mem.mem_outb[0] = 1'b0;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_20.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_40.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_42.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_64.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_74.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_112.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_114.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_top_track_122.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_26.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_38.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_42.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_52.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_60.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_62.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_76.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_84.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_90.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_92.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_98.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_100.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__0_.mem_right_track_102.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_106.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_108.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_110.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_112.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_128.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_132.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_138.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_140.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__1_.mem_top_track_8.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__1_.mem_top_track_16.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_24.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_0__1_.mem_top_track_32.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__1_.mem_top_track_40.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__1_.mem_top_track_48.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_56.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_64.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__1_.mem_top_track_72.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.sb_0__1_.mem_top_track_80.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__1_.mem_top_track_88.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_0__1_.mem_top_track_96.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_top_track_104.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__1_.mem_top_track_112.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_0__1_.mem_top_track_120.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__1_.mem_top_track_128.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__1_.mem_top_track_136.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_0__1_.mem_top_track_144.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__1_.mem_right_track_58.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_60.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_66.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_74.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_78.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_84.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_90.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_92.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_94.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_96.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_98.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_100.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_108.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__1_.mem_right_track_114.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_116.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_122.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_124.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__1_.mem_right_track_126.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_132.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__1_.mem_right_track_138.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_25.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_41.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_97.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__2_.mem_top_track_24.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_42.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_58.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_60.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_66.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__2_.mem_right_track_68.mem_outb[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_74.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_84.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_90.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_94.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_98.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_100.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_104.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__2_.mem_right_track_106.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_108.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_114.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_122.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_124.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_132.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_134.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_136.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_138.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_0__2_.mem_right_track_144.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_top_track_40.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_top_track_104.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_58.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_68.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_74.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_80.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_84.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_88.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_98.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_102.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_106.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_108.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_114.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__3_.mem_right_track_122.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_124.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_128.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_9.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_17.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_25.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_49.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_57.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_65.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_81.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_105.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_121.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_129.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_0__4_.mem_top_track_56.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_58.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_60.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_64.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_66.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_74.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_84.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__4_.mem_right_track_90.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_94.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_98.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_100.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_102.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_108.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_112.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_114.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_122.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_124.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_132.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_138.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_0__4_.mem_right_track_140.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_41.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_57.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_65.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_97.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_105.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_113.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_121.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_42.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_58.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_60.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_62.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_66.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_68.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_70.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_74.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_76.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_78.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_82.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_84.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_86.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_90.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_92.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_94.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_98.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_100.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_102.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_106.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_108.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_110.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_114.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_116.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_118.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_122.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_124.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_126.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_130.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_132.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_134.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_136.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_0__5_.mem_right_track_138.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_140.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_142.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_33.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_41.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_113.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_121.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_137.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_42.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_66.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_80.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_108.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_130.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_right_track_138.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_right_track_140.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_144.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_77.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_77.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_85.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_85.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_105.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_107.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_107.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_111.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_111.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_133.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_133.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_137.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_0__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_64.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_82.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_98.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_100.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_120.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_122.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_132.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__0_.mem_top_track_138.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_16.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_32.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_64.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_88.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__0_.mem_right_track_96.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__0_.mem_right_track_112.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__0_.mem_right_track_128.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_8.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_24.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_40.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_top_track_48.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_top_track_64.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__1_.mem_top_track_72.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_80.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_1__1_.mem_top_track_88.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_top_track_96.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__1_.mem_top_track_104.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_top_track_112.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__1_.mem_top_track_120.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_1__1_.mem_top_track_128.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__1_.mem_top_track_136.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_1__1_.mem_top_track_144.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_8.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_right_track_72.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__1_.mem_right_track_112.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_17.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_25.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_33.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_41.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_129.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__1_.mem_bottom_track_145.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_1__1_.mem_left_track_9.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__1_.mem_left_track_17.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_left_track_25.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__1_.mem_left_track_33.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_41.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_left_track_49.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__1_.mem_left_track_65.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_left_track_73.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__1_.mem_left_track_81.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__1_.mem_left_track_129.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__1_.mem_left_track_137.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__1_.mem_left_track_145.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__2_.mem_top_track_8.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__2_.mem_top_track_16.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__2_.mem_top_track_24.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__2_.mem_top_track_40.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__2_.mem_top_track_120.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__2_.mem_right_track_8.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__2_.mem_right_track_32.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__2_.mem_right_track_48.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__2_.mem_right_track_64.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__2_.mem_right_track_88.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__2_.mem_right_track_96.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__2_.mem_right_track_112.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__2_.mem_right_track_136.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_17.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__2_.mem_left_track_17.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__2_.mem_left_track_25.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__2_.mem_left_track_49.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_left_track_73.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_81.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_left_track_113.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_121.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.sb_1__2_.mem_left_track_137.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__2_.mem_left_track_145.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_top_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__3_.mem_top_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__3_.mem_right_track_8.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_16.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_24.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_64.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__3_.mem_right_track_88.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_right_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__3_.mem_right_track_136.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_17.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_25.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_33.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_57.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_65.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_73.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_89.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_137.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_1__3_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_left_track_97.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_left_track_129.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__3_.mem_left_track_145.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__4_.mem_right_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_right_track_104.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_1__4_.mem_right_track_136.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_9.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_25.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_33.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_81.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_97.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.sb_1__4_.mem_left_track_97.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__4_.mem_left_track_121.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_1__5_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__5_.mem_right_track_144.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_33.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_41.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_65.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_81.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_89.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_105.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_121.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_129.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_1__5_.mem_left_track_9.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_1__6_.mem_right_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_1__6_.mem_right_track_40.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_9.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_49.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_59.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_59.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_1__6_.mem_bottom_track_145.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_1__6_.mem_left_track_41.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_74.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_86.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_90.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_98.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_98.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_100.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_114.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_122.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_124.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_128.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_134.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__0_.mem_top_track_136.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_16.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_56.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_72.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_right_track_88.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_96.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_right_track_120.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_right_track_128.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_right_track_144.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_left_track_9.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_33.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_41.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_left_track_65.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_left_track_73.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_89.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__0_.mem_left_track_97.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_left_track_105.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__0_.mem_left_track_113.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__0_.mem_left_track_129.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__1_.mem_top_track_16.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__1_.mem_top_track_24.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_32.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_48.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_top_track_64.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_72.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_top_track_80.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_top_track_88.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_top_track_104.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_top_track_112.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__1_.mem_top_track_120.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__1_.mem_top_track_136.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_top_track_144.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_8.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_40.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_80.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_right_track_96.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_right_track_112.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_right_track_120.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_17.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_25.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_41.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_137.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_bottom_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__1_.mem_left_track_9.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__1_.mem_left_track_17.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__1_.mem_left_track_41.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__1_.mem_left_track_49.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__1_.mem_left_track_57.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_left_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__1_.mem_left_track_89.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__1_.mem_left_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__1_.mem_left_track_121.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__1_.mem_left_track_129.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__1_.mem_left_track_137.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__1_.mem_left_track_145.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_top_track_16.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_top_track_24.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_top_track_40.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_top_track_48.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_top_track_64.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__2_.mem_top_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_top_track_112.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_top_track_120.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_top_track_128.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_top_track_136.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_24.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_right_track_48.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_64.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_right_track_88.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_right_track_144.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_9.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_17.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_33.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_41.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_57.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_65.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_105.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_113.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_137.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_left_track_17.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__2_.mem_left_track_25.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_left_track_49.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_left_track_65.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_left_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__2_.mem_left_track_81.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__2_.mem_left_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__2_.mem_left_track_113.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__2_.mem_left_track_129.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__2_.mem_left_track_137.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_top_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__3_.mem_right_track_40.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_64.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_right_track_80.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_right_track_112.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_right_track_120.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__3_.mem_right_track_136.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_9.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_89.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_129.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_137.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_bottom_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_9.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_left_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__3_.mem_left_track_65.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__3_.mem_left_track_89.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__4_.mem_top_track_16.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_top_track_48.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_right_track_8.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_right_track_16.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_24.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__4_.mem_right_track_40.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__4_.mem_right_track_80.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_right_track_96.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__4_.mem_right_track_120.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_49.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_73.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_81.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_97.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_105.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__4_.mem_left_track_33.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_2__4_.mem_left_track_121.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__4_.mem_left_track_137.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_right_track_24.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_right_track_56.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_right_track_72.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_80.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_104.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_right_track_112.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_128.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_17.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_73.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_89.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_137.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_2__5_.mem_left_track_57.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_2__5_.mem_left_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__6_.mem_right_track_8.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_2__6_.mem_right_track_72.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_33.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_43.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_43.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_99.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_99.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_105.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_2__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_2__6_.mem_left_track_25.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__6_.mem_left_track_49.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_2__6_.mem_left_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_54.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_56.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_60.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_66.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_68.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_72.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_74.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_88.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_90.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_92.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_96.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_96.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_112.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_120.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_122.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__0_.mem_top_track_124.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_126.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_130.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_16.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_24.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_40.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_right_track_72.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_88.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_96.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_112.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_120.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_right_track_128.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_right_track_144.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_left_track_9.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_17.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_25.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_left_track_33.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_left_track_41.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_3__0_.mem_left_track_57.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__0_.mem_left_track_73.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_left_track_105.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_113.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_121.mem_outb[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__0_.mem_left_track_137.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__1_.mem_top_track_8.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_3__1_.mem_top_track_16.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__1_.mem_top_track_24.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__1_.mem_top_track_32.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__1_.mem_top_track_40.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__1_.mem_top_track_48.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_3__1_.mem_top_track_56.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__1_.mem_top_track_64.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_3__1_.mem_top_track_72.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__1_.mem_top_track_80.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__1_.mem_top_track_88.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__1_.mem_top_track_96.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__1_.mem_top_track_104.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__1_.mem_top_track_112.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_top_track_120.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__1_.mem_top_track_128.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_3__1_.mem_top_track_136.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__1_.mem_top_track_144.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_8.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.sb_3__1_.mem_right_track_24.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__1_.mem_right_track_72.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_80.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_88.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_104.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_120.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__1_.mem_right_track_128.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_3__1_.mem_right_track_136.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__1_.mem_right_track_144.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_9.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_73.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_105.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_113.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_bottom_track_145.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_left_track_9.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__1_.mem_left_track_17.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_3__1_.mem_left_track_25.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_left_track_41.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__1_.mem_left_track_49.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__1_.mem_left_track_65.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__1_.mem_left_track_81.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_105.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__1_.mem_left_track_121.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__1_.mem_left_track_137.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_top_track_8.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__2_.mem_top_track_24.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_3__2_.mem_top_track_72.mem_outb[0:3] = 4'b1010;
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__2_.mem_top_track_88.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__2_.mem_top_track_96.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__2_.mem_top_track_120.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__2_.mem_top_track_136.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_top_track_144.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__2_.mem_right_track_16.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_right_track_40.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__2_.mem_right_track_48.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_right_track_96.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_right_track_104.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_128.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_17.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_121.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__2_.mem_left_track_17.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__2_.mem_left_track_25.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__2_.mem_left_track_33.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__2_.mem_left_track_41.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_left_track_65.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__2_.mem_left_track_73.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__2_.mem_left_track_97.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__2_.mem_left_track_105.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_left_track_113.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__2_.mem_left_track_121.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__2_.mem_left_track_129.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_3__2_.mem_left_track_137.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__3_.mem_top_track_8.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_top_track_56.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_3__3_.mem_top_track_80.mem_outb[0:3] = 4'b1100;
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_16.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_24.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_right_track_32.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_right_track_56.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_right_track_88.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_120.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_right_track_128.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_3__3_.mem_right_track_144.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_25.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_49.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_89.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_97.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_105.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_121.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_left_track_9.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_3__3_.mem_left_track_25.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_left_track_49.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__3_.mem_left_track_73.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__3_.mem_left_track_129.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_3__4_.mem_top_track_112.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__4_.mem_right_track_40.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_72.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__4_.mem_right_track_104.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__4_.mem_right_track_144.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_9.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_73.mem_outb[0:3] = 4'b0100;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_81.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_89.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_105.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_113.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_3__4_.mem_left_track_25.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_3__4_.mem_left_track_73.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_3__4_.mem_left_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_8.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_32.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_40.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_48.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_56.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_64.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_72.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_80.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_88.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_96.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_104.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_112.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_144.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_3__5_.mem_right_track_8.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__5_.mem_right_track_40.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_3__5_.mem_right_track_48.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_3__5_.mem_right_track_104.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_120.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_17.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_97.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_105.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_113.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_137.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_145.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_3__5_.mem_left_track_81.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_3__6_.mem_right_track_88.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_9.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_3__6_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_35.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_113.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_121.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_38.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_52.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_56.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_60.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_62.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_64.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_66.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_68.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_70.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_74.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_76.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_78.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_80.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_82.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_84.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_86.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_88.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_92.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_94.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_96.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_98.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_100.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_102.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_104.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_106.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_110.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_112.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_114.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_116.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_118.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_120.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_122.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_124.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_128.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__0_.mem_top_track_130.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_132.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_134.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_136.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_138.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_140.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_142.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_9.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_17.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_19.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_19.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_27.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_27.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_33.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_35.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_35.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_49.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_53.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_65.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_73.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_89.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_97.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_105.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_107.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_107.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_113.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_121.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_123.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_123.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_129.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_131.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_131.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_137.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_4__1_.mem_top_track_8.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_4__1_.mem_top_track_16.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_4__1_.mem_top_track_24.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__1_.mem_top_track_32.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.sb_4__1_.mem_top_track_40.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_4__1_.mem_top_track_48.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__1_.mem_top_track_56.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__1_.mem_top_track_64.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__1_.mem_top_track_72.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.sb_4__1_.mem_top_track_80.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__1_.mem_top_track_88.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_4__1_.mem_top_track_96.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_4__1_.mem_top_track_104.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__1_.mem_top_track_112.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_4__1_.mem_top_track_120.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_4__1_.mem_top_track_128.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_4__1_.mem_top_track_136.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_4__1_.mem_top_track_144.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_17.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_25.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_49.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_65.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_105.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_113.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_121.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_129.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__1_.mem_bottom_track_145.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_3.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_3.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_5.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__1_.mem_left_track_5.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_9.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_11.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_11.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_15.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_15.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_17.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_19.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_19.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_21.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__1_.mem_left_track_21.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__1_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_27.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__1_.mem_left_track_27.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_31.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_31.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_37.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_37.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_39.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_39.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_41.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_43.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_43.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_53.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_53.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_57.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_59.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_59.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_61.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_61.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_65.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_69.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_69.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_75.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_left_track_75.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_81.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_83.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_83.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_93.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_93.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__1_.mem_left_track_97.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__1_.mem_left_track_99.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_99.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_103.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__1_.mem_left_track_103.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_107.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_107.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__1_.mem_left_track_113.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__1_.mem_left_track_115.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__1_.mem_left_track_115.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__1_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__1_.mem_left_track_121.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__1_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_127.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__1_.mem_left_track_127.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_131.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__1_.mem_left_track_131.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__1_.mem_left_track_133.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_133.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__1_.mem_left_track_137.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__1_.mem_left_track_139.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__1_.mem_left_track_139.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__1_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__1_.mem_left_track_145.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__2_.mem_top_track_40.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__2_.mem_top_track_48.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__2_.mem_top_track_72.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__2_.mem_top_track_88.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__2_.mem_top_track_128.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__2_.mem_top_track_136.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__2_.mem_top_track_144.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_9.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_17.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_25.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_33.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_41.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_49.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_57.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_65.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_73.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_81.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_89.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_97.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_105.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_113.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_121.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_129.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_137.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__2_.mem_bottom_track_145.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_3.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_left_track_3.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_7.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_7.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_19.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_19.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_27.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_left_track_27.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_35.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_35.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_39.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__2_.mem_left_track_39.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_43.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_43.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_left_track_49.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_left_track_51.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_51.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_53.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_53.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_57.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_59.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__2_.mem_left_track_59.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__2_.mem_left_track_61.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_61.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_left_track_65.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_69.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__2_.mem_left_track_69.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__2_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_75.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_75.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_77.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_77.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_out[0:3] = 4'b1010;
	force U0_formal_verification.sb_4__2_.mem_left_track_81.mem_outb[0:3] = 4'b0101;
	force U0_formal_verification.sb_4__2_.mem_left_track_83.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_83.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_85.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__2_.mem_left_track_85.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__2_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_91.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_91.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_99.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__2_.mem_left_track_99.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__2_.mem_left_track_101.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_left_track_101.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_105.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_107.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_107.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__2_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_113.mem_outb[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_125.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_4__2_.mem_left_track_125.mem_outb[0:3] = 4'b0110;
	force U0_formal_verification.sb_4__2_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_left_track_129.mem_outb[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_left_track_131.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.sb_4__2_.mem_left_track_131.mem_outb[0:3] = 4'b1101;
	force U0_formal_verification.sb_4__2_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_135.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.sb_4__2_.mem_left_track_135.mem_outb[0:3] = 4'b0001;
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_139.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_139.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.sb_4__2_.mem_left_track_145.mem_outb[0:3] = 4'b1011;
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_top_track_32.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_top_track_72.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_top_track_80.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_96.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_top_track_112.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_128.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_9.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_25.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_33.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_41.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_out[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_49.mem_outb[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_57.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_65.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_73.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_81.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_89.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_97.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_105.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_113.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_121.mem_outb[0:2] = 3'b100;
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_129.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_5.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_11.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_17.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_23.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_23.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_35.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_35.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_41.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_53.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_53.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_71.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_71.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_83.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_83.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_89.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_95.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_95.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_105.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_107.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__3_.mem_left_track_107.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__3_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_125.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_125.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_143.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_143.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_96.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_104.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_112.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__4_.mem_top_track_120.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_128.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_136.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_144.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_9.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_17.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_25.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_33.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_41.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_49.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_57.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_65.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_73.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_81.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_89.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_97.mem_outb[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_105.mem_outb[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_113.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_121.mem_outb[0:2] = 3'b101;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_129.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_137.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_145.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_27.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_27.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_35.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_35.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_67.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__4_.mem_left_track_67.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__4_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__4_.mem_left_track_73.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__4_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_91.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__4_.mem_left_track_91.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__4_.mem_left_track_93.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_93.mem_outb[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_8.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_16.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_24.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_32.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_40.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_48.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_56.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_64.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_72.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_80.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_88.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__5_.mem_top_track_96.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_104.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_112.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_120.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_4__5_.mem_top_track_128.mem_outb[0:2] = 3'b110;
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_136.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_144.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_25.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_33.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_73.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_81.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_97.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_105.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_113.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_121.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_129.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_137.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.sb_4__5_.mem_bottom_track_145.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_3.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_5.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_7.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_9.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_11.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_13.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_15.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_17.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_19.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_19.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_21.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_23.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_23.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_25.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_27.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__5_.mem_left_track_27.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_29.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_31.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_31.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_33.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_35.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_4__5_.mem_left_track_35.mem_outb[0:3] = 4'b1000;
	force U0_formal_verification.sb_4__5_.mem_left_track_37.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_37.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_39.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_39.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_41.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_43.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_43.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_45.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_45.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_47.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_47.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_49.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_51.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_51.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_53.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_53.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_55.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_55.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_57.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_59.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_59.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_61.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_61.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_63.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_63.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_65.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_67.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_67.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_69.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_69.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_71.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_71.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_73.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_75.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_75.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_77.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_77.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_79.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_79.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_81.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_83.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_83.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_85.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_85.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_87.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_87.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_89.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_91.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_91.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_93.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_93.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_95.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_95.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_97.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_99.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_99.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_101.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_101.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_103.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_103.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_105.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_107.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_107.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_109.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_109.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_111.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_111.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_113.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_115.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_115.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_117.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_117.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_119.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_119.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_121.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_123.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_123.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_125.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_125.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_127.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_127.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_129.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_131.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_131.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_133.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_133.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_135.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_135.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_137.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_139.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_139.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_141.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_141.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_143.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_143.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_145.mem_outb[0:3] = {4{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_9.mem_outb[0:1] = 2'b01;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_11.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_43.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_43.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_73.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_87.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_87.mem_outb[0:1] = 2'b10;
	force U0_formal_verification.sb_4__6_.mem_bottom_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_3.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_5.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_5.mem_outb[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_7.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_9.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_11.mem_outb[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_13.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_15.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_17.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_19.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_21.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_23.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_25.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_27.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_29.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_31.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_33.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_37.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_39.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_41.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_43.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_45.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_47.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_49.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_51.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_55.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_57.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_59.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_61.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_61.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_63.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_63.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_65.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_67.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_67.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_69.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_69.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_73.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_75.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_75.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_77.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_77.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_79.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_79.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_81.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_83.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_83.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_85.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_85.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_87.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_87.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_91.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_91.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_93.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_93.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_95.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_95.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_97.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_99.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_99.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_101.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_101.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_103.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_103.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_105.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_109.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_109.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_111.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_111.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_113.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_115.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_115.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_117.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_117.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_119.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_119.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_121.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_123.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_123.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_127.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_127.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_129.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_131.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_131.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_133.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_133.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_135.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_135.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_137.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_139.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_139.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_141.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_141.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_145.mem_outb[0:1] = {2{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_0.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_1.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_19.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_19.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_20.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_20.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_21.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_21.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_22.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_22.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_23.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_23.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_24.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_24.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_25.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_25.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_26.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_26.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_27.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_27.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_28.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_28.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_29.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_29.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_30.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_30.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_31.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_31.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_32.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_32.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_33.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_33.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_34.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_34.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_35.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_35.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_70.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_70.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_71.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_71.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_72.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_72.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_73.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_73.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_74.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_74.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_75.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_75.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_76.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_76.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_77.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_77.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_78.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_78.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_79.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_79.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_80.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_80.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_81.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_81.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_82.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_82.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_83.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_83.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_84.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_84.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_85.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_85.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_86.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_86.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_bottom_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_19.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_19.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_20.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_20.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_21.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_21.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_22.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_22.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_23.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_23.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_24.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_24.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_25.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_25.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_26.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_26.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_27.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_27.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_28.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_28.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_29.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_29.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_30.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_30.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_31.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_31.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_32.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_32.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_33.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_33.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_34.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_34.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_35.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_35.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_70.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_70.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_71.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_71.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_72.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_72.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_73.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_73.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_74.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_74.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_75.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_75.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_76.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_76.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_77.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_77.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_78.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_78.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_79.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_79.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_80.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_80.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_81.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_81.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_82.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_82.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_83.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_83.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_84.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_84.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_85.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_85.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_86.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_86.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_bottom_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_4.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_6.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_7.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cbx_3__0_.mem_bottom_ipin_1.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_4.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_5.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_6.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_7.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_4.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_5.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_6.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_7.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_0.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_1.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_53.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_53.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_54.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_54.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_55.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_55.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_56.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_56.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_57.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_57.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_58.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_58.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_59.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_59.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_60.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_60.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_61.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_61.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_62.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_62.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_63.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_63.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_64.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_64.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_65.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_65.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_66.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_66.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_67.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_67.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_68.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_68.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_69.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_69.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_bottom_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_53.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_53.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_54.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_54.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_55.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_55.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_56.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_56.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_57.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_57.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_58.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_58.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_59.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_59.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_60.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_60.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_61.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_61.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_62.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_62.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_63.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_63.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_64.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_64.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_65.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_65.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_66.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_66.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_67.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_67.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_68.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_68.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_69.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_69.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_bottom_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_89.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_89.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_bottom_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_0.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_18.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_18.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_19.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_19.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_20.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_20.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_21.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_21.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_22.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_22.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_23.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_23.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_24.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_24.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_25.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_25.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_26.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_26.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_27.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_27.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_28.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_28.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_29.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_29.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_30.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_30.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_31.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_31.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_32.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_32.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_33.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_33.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_34.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_34.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_69.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_69.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_70.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_70.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_71.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_71.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_72.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_72.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_73.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_73.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_74.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_74.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_75.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_75.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_76.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_76.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_77.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_77.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_78.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_78.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_79.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_79.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_80.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_80.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_81.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_81.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_82.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_82.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_83.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_83.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_84.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_84.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_85.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_85.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_0__2_.mem_left_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_left_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_left_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_19.mem_out[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_19.mem_outb[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_20.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_20.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_21.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_21.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_22.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_22.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_23.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_23.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_24.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_24.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_25.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_25.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_26.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_26.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_27.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_27.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_28.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_28.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_29.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_29.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_30.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_30.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_31.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_31.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_32.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_32.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_33.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_33.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_34.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_34.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_35.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_35.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_70.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_70.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_71.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_71.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_72.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_72.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_73.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_73.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_74.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_74.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_75.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_75.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_76.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_76.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_77.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_77.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_78.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_78.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_79.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_79.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_80.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_80.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_81.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_81.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_82.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_82.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_83.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_83.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_84.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_84.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_85.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_85.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_86.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_86.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cby_1__2_.mem_right_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_0.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_52.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_52.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_53.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_53.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_54.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_54.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_55.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_55.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_56.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_56.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_57.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_57.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_58.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_58.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_59.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_59.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_60.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_60.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_61.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_61.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_62.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_62.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_63.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_63.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_64.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_64.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_65.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_65.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_66.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_66.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_67.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_67.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_68.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_68.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_3__2_.mem_left_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_left_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_left_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_left_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_0.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_1.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_out[0:4] = 5'b00101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_2.mem_outb[0:4] = 5'b11010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_3.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_4.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_5.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_6.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__1_.mem_left_ipin_7.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_out[0:4] = 5'b10110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_0.mem_outb[0:4] = 5'b01001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_1.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_2.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_3.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_4.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_5.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_6.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__2_.mem_left_ipin_7.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_53.mem_out[0:4] = 5'b01111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_53.mem_outb[0:4] = 5'b10000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_54.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_54.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_55.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_55.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_56.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_56.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_57.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_57.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_58.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_58.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_59.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_59.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_60.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_60.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_61.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_61.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_62.mem_out[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_62.mem_outb[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_63.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_63.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_64.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_64.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_65.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_65.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_66.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_66.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_67.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_67.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_68.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_68.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_69.mem_out[0:4] = 5'b01001;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_69.mem_outb[0:4] = 5'b10110;
	force U0_formal_verification.cby_4__2_.mem_right_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_0.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_out[0:4] = 5'b01011;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_1.mem_outb[0:4] = 5'b10100;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_2.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_2.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_3.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_3.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_4.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_4.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_5.mem_out[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_5.mem_outb[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_6.mem_out[0:4] = 5'b00100;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_6.mem_outb[0:4] = 5'b11011;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_7.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__3_.mem_left_ipin_7.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_0.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_out[0:4] = 5'b00111;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_1.mem_outb[0:4] = 5'b11000;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_2.mem_out[0:4] = 5'b11010;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_2.mem_outb[0:4] = 5'b00101;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_3.mem_out[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_3.mem_outb[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_4.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_4.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_5.mem_out[0:4] = 5'b00011;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_5.mem_outb[0:4] = 5'b11100;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_6.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_6.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_7.mem_out[0:4] = 5'b11001;
	force U0_formal_verification.cby_4__4_.mem_left_ipin_7.mem_outb[0:4] = 5'b00110;
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_0.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_out[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_1.mem_outb[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_2.mem_out[0:4] = 5'b10101;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_2.mem_outb[0:4] = 5'b01010;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_3.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_3.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_4.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_4.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_5.mem_out[0:4] = 5'b10011;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_5.mem_outb[0:4] = 5'b01100;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_6.mem_out[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_6.mem_outb[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_7.mem_out[0:4] = 5'b11011;
	force U0_formal_verification.cby_4__5_.mem_left_ipin_7.mem_outb[0:4] = 5'b00100;
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_16.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_16.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_17.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_17.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_18.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_18.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_19.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_19.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_20.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_20.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_21.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_21.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_22.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_22.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_23.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_23.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_24.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_24.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_25.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_25.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_26.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_26.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_27.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_27.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_28.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_28.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_29.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_29.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_30.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_30.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_31.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_31.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_32.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_32.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_33.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_33.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_34.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_34.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_35.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_35.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_36.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_36.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_37.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_37.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_38.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_38.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_39.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_39.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_40.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_40.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_41.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_41.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_42.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_42.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_43.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_43.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_44.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_44.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_45.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_45.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_46.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_46.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_47.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_47.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_48.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_48.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_49.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_49.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_50.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_50.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_51.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_51.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_52.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_52.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_53.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_53.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_54.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_54.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_55.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_55.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_56.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_56.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_57.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_57.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_58.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_58.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_59.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_59.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_60.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_60.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_61.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_61.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_62.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_62.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_63.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_63.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_64.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_64.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_65.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_65.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_66.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_66.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_67.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_67.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_68.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_68.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_69.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_69.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_70.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_70.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_71.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_71.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_72.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_72.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_73.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_73.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_74.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_74.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_75.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_75.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_76.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_76.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_77.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_77.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_78.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_78.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_79.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_79.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_80.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_80.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_81.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_81.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_82.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_82.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_83.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_83.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_84.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_84.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_85.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_85.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_86.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_86.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_87.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_87.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_88.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_88.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_out[0:4] = 5'b11110;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_0.mem_outb[0:4] = 5'b00001;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_out[0:4] = 5'b01110;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_1.mem_outb[0:4] = 5'b10001;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_2.mem_out[0:4] = 5'b10111;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_2.mem_outb[0:4] = 5'b01000;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_3.mem_out[0:4] = 5'b01101;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_3.mem_outb[0:4] = 5'b10010;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_4.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_4.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_5.mem_out[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_5.mem_outb[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_6.mem_out[0:4] = 5'b10001;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_6.mem_outb[0:4] = 5'b01110;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_7.mem_out[0:4] = 5'b00010;
	force U0_formal_verification.cby_4__6_.mem_left_ipin_7.mem_outb[0:4] = 5'b11101;
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_outb[0:4] = {5{1'b1}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:4] = {5{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_outb[0:4] = {5{1'b1}};
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for router_tb_top_formal_verification -----

//----- Default net type -----
`default_nettype wire

