//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for pb_type: router_wrap_slice
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sun Jul 21 19:29:39 2024
//-------------------------------------------
// ----- BEGIN Physical programmable logic block Verilog module: router_wrap_slice -----
//----- Default net type -----
`default_nettype none

// ----- Verilog module for logical_tile_router_mode_router_wrap__router_wrap_slice -----
module logical_tile_router_mode_router_wrap__router_wrap_slice(clk,
                                                               set,
                                                               reset,
                                                               prog_clk,
                                                               router_wrap_slice_RST__cfg,
                                                               router_wrap_slice_MY_XPOS_cfg,
                                                               router_wrap_slice_MY_YPOS_cfg,
                                                               router_wrap_slice_IDATA_0_cfg,
                                                               router_wrap_slice_IDATA_1_cfg,
                                                               router_wrap_slice_IDATA_2_cfg,
                                                               router_wrap_slice_IDATA_3_cfg,
                                                               router_wrap_slice_IDATA_4_cfg,
                                                               router_wrap_slice_IVALID_0_cfg,
                                                               router_wrap_slice_IVALID_1_cfg,
                                                               router_wrap_slice_IVALID_2_cfg,
                                                               router_wrap_slice_IVALID_3_cfg,
                                                               router_wrap_slice_IVALID_4_cfg,
                                                               router_wrap_slice_IVCH_0_cfg,
                                                               router_wrap_slice_IVCH_1_cfg,
                                                               router_wrap_slice_IVCH_2_cfg,
                                                               router_wrap_slice_IVCH_3_cfg,
                                                               router_wrap_slice_IVCH_4_cfg,
                                                               router_wrap_slice_IACK_0_cfg,
                                                               router_wrap_slice_IACK_1_cfg,
                                                               router_wrap_slice_IACK_2_cfg,
                                                               router_wrap_slice_IACK_3_cfg,
                                                               router_wrap_slice_IACK_4_cfg,
                                                               router_wrap_slice_ILCK_0_cfg,
                                                               router_wrap_slice_ILCK_1_cfg,
                                                               router_wrap_slice_ILCK_2_cfg,
                                                               router_wrap_slice_ILCK_3_cfg,
                                                               router_wrap_slice_ILCK_4_cfg,
                                                               router_wrap_slice_clk,
                                                               ccff_head,
                                                               router_wrap_slice_ODATA_0_cfg,
                                                               router_wrap_slice_ODATA_1_cfg,
                                                               router_wrap_slice_ODATA_2_cfg,
                                                               router_wrap_slice_ODATA_3_cfg,
                                                               router_wrap_slice_ODATA_4_cfg,
                                                               router_wrap_slice_OVALID_0_cfg,
                                                               router_wrap_slice_OVALID_1_cfg,
                                                               router_wrap_slice_OVALID_2_cfg,
                                                               router_wrap_slice_OVALID_3_cfg,
                                                               router_wrap_slice_OVALID_4_cfg,
                                                               router_wrap_slice_OVCH_0_cfg,
                                                               router_wrap_slice_OVCH_1_cfg,
                                                               router_wrap_slice_OVCH_2_cfg,
                                                               router_wrap_slice_OVCH_3_cfg,
                                                               router_wrap_slice_OVCH_4_cfg,
                                                               router_wrap_slice_OACK_0_cfg,
                                                               router_wrap_slice_OACK_1_cfg,
                                                               router_wrap_slice_OACK_2_cfg,
                                                               router_wrap_slice_OACK_3_cfg,
                                                               router_wrap_slice_OACK_4_cfg,
                                                               router_wrap_slice_ORDY_0_cfg,
                                                               router_wrap_slice_ORDY_1_cfg,
                                                               router_wrap_slice_ORDY_2_cfg,
                                                               router_wrap_slice_ORDY_3_cfg,
                                                               router_wrap_slice_ORDY_4_cfg,
                                                               router_wrap_slice_OLCK_0_cfg,
                                                               router_wrap_slice_OLCK_1_cfg,
                                                               router_wrap_slice_OLCK_2_cfg,
                                                               router_wrap_slice_OLCK_3_cfg,
                                                               router_wrap_slice_OLCK_4_cfg,
                                                               ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] set;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_RST__cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_MY_XPOS_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_MY_YPOS_cfg;
//----- INPUT PORTS -----
input [0:34] router_wrap_slice_IDATA_0_cfg;
//----- INPUT PORTS -----
input [0:34] router_wrap_slice_IDATA_1_cfg;
//----- INPUT PORTS -----
input [0:34] router_wrap_slice_IDATA_2_cfg;
//----- INPUT PORTS -----
input [0:34] router_wrap_slice_IDATA_3_cfg;
//----- INPUT PORTS -----
input [0:34] router_wrap_slice_IDATA_4_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVALID_0_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVALID_1_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVALID_2_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVALID_3_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVALID_4_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVCH_0_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVCH_1_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVCH_2_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVCH_3_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_IVCH_4_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_IACK_0_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_IACK_1_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_IACK_2_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_IACK_3_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_IACK_4_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_ILCK_0_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_ILCK_1_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_ILCK_2_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_ILCK_3_cfg;
//----- INPUT PORTS -----
input [0:1] router_wrap_slice_ILCK_4_cfg;
//----- INPUT PORTS -----
input [0:0] router_wrap_slice_clk;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:34] router_wrap_slice_ODATA_0_cfg;
//----- OUTPUT PORTS -----
output [0:34] router_wrap_slice_ODATA_1_cfg;
//----- OUTPUT PORTS -----
output [0:34] router_wrap_slice_ODATA_2_cfg;
//----- OUTPUT PORTS -----
output [0:34] router_wrap_slice_ODATA_3_cfg;
//----- OUTPUT PORTS -----
output [0:34] router_wrap_slice_ODATA_4_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVALID_0_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVALID_1_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVALID_2_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVALID_3_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVALID_4_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVCH_0_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVCH_1_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVCH_2_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVCH_3_cfg;
//----- OUTPUT PORTS -----
output [0:0] router_wrap_slice_OVCH_4_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OACK_0_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OACK_1_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OACK_2_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OACK_3_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OACK_4_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_ORDY_0_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_ORDY_1_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_ORDY_2_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_ORDY_3_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_ORDY_4_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OLCK_0_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OLCK_1_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OLCK_2_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OLCK_3_cfg;
//----- OUTPUT PORTS -----
output [0:1] router_wrap_slice_OLCK_4_cfg;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
wire [0:0] router_wrap_slice_RST__cfg;
wire [0:1] router_wrap_slice_MY_XPOS_cfg;
wire [0:1] router_wrap_slice_MY_YPOS_cfg;
wire [0:34] router_wrap_slice_IDATA_0_cfg;
wire [0:34] router_wrap_slice_IDATA_1_cfg;
wire [0:34] router_wrap_slice_IDATA_2_cfg;
wire [0:34] router_wrap_slice_IDATA_3_cfg;
wire [0:34] router_wrap_slice_IDATA_4_cfg;
wire [0:0] router_wrap_slice_IVALID_0_cfg;
wire [0:0] router_wrap_slice_IVALID_1_cfg;
wire [0:0] router_wrap_slice_IVALID_2_cfg;
wire [0:0] router_wrap_slice_IVALID_3_cfg;
wire [0:0] router_wrap_slice_IVALID_4_cfg;
wire [0:0] router_wrap_slice_IVCH_0_cfg;
wire [0:0] router_wrap_slice_IVCH_1_cfg;
wire [0:0] router_wrap_slice_IVCH_2_cfg;
wire [0:0] router_wrap_slice_IVCH_3_cfg;
wire [0:0] router_wrap_slice_IVCH_4_cfg;
wire [0:1] router_wrap_slice_IACK_0_cfg;
wire [0:1] router_wrap_slice_IACK_1_cfg;
wire [0:1] router_wrap_slice_IACK_2_cfg;
wire [0:1] router_wrap_slice_IACK_3_cfg;
wire [0:1] router_wrap_slice_IACK_4_cfg;
wire [0:1] router_wrap_slice_ILCK_0_cfg;
wire [0:1] router_wrap_slice_ILCK_1_cfg;
wire [0:1] router_wrap_slice_ILCK_2_cfg;
wire [0:1] router_wrap_slice_ILCK_3_cfg;
wire [0:1] router_wrap_slice_ILCK_4_cfg;
wire [0:0] router_wrap_slice_clk;
wire [0:34] router_wrap_slice_ODATA_0_cfg;
wire [0:34] router_wrap_slice_ODATA_1_cfg;
wire [0:34] router_wrap_slice_ODATA_2_cfg;
wire [0:34] router_wrap_slice_ODATA_3_cfg;
wire [0:34] router_wrap_slice_ODATA_4_cfg;
wire [0:0] router_wrap_slice_OVALID_0_cfg;
wire [0:0] router_wrap_slice_OVALID_1_cfg;
wire [0:0] router_wrap_slice_OVALID_2_cfg;
wire [0:0] router_wrap_slice_OVALID_3_cfg;
wire [0:0] router_wrap_slice_OVALID_4_cfg;
wire [0:0] router_wrap_slice_OVCH_0_cfg;
wire [0:0] router_wrap_slice_OVCH_1_cfg;
wire [0:0] router_wrap_slice_OVCH_2_cfg;
wire [0:0] router_wrap_slice_OVCH_3_cfg;
wire [0:0] router_wrap_slice_OVCH_4_cfg;
wire [0:1] router_wrap_slice_OACK_0_cfg;
wire [0:1] router_wrap_slice_OACK_1_cfg;
wire [0:1] router_wrap_slice_OACK_2_cfg;
wire [0:1] router_wrap_slice_OACK_3_cfg;
wire [0:1] router_wrap_slice_OACK_4_cfg;
wire [0:1] router_wrap_slice_ORDY_0_cfg;
wire [0:1] router_wrap_slice_ORDY_1_cfg;
wire [0:1] router_wrap_slice_ORDY_2_cfg;
wire [0:1] router_wrap_slice_ORDY_3_cfg;
wire [0:1] router_wrap_slice_ORDY_4_cfg;
wire [0:1] router_wrap_slice_OLCK_0_cfg;
wire [0:1] router_wrap_slice_OLCK_1_cfg;
wire [0:1] router_wrap_slice_OLCK_2_cfg;
wire [0:1] router_wrap_slice_OLCK_3_cfg;
wire [0:1] router_wrap_slice_OLCK_4_cfg;
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:0] direct_interc_0_out;
wire [0:0] direct_interc_100_out;
wire [0:0] direct_interc_101_out;
wire [0:0] direct_interc_102_out;
wire [0:0] direct_interc_103_out;
wire [0:0] direct_interc_104_out;
wire [0:0] direct_interc_105_out;
wire [0:0] direct_interc_106_out;
wire [0:0] direct_interc_107_out;
wire [0:0] direct_interc_108_out;
wire [0:0] direct_interc_109_out;
wire [0:0] direct_interc_10_out;
wire [0:0] direct_interc_110_out;
wire [0:0] direct_interc_111_out;
wire [0:0] direct_interc_112_out;
wire [0:0] direct_interc_113_out;
wire [0:0] direct_interc_114_out;
wire [0:0] direct_interc_115_out;
wire [0:0] direct_interc_116_out;
wire [0:0] direct_interc_117_out;
wire [0:0] direct_interc_118_out;
wire [0:0] direct_interc_119_out;
wire [0:0] direct_interc_11_out;
wire [0:0] direct_interc_120_out;
wire [0:0] direct_interc_121_out;
wire [0:0] direct_interc_122_out;
wire [0:0] direct_interc_123_out;
wire [0:0] direct_interc_124_out;
wire [0:0] direct_interc_125_out;
wire [0:0] direct_interc_126_out;
wire [0:0] direct_interc_127_out;
wire [0:0] direct_interc_128_out;
wire [0:0] direct_interc_129_out;
wire [0:0] direct_interc_12_out;
wire [0:0] direct_interc_130_out;
wire [0:0] direct_interc_131_out;
wire [0:0] direct_interc_132_out;
wire [0:0] direct_interc_133_out;
wire [0:0] direct_interc_134_out;
wire [0:0] direct_interc_135_out;
wire [0:0] direct_interc_136_out;
wire [0:0] direct_interc_137_out;
wire [0:0] direct_interc_138_out;
wire [0:0] direct_interc_139_out;
wire [0:0] direct_interc_13_out;
wire [0:0] direct_interc_140_out;
wire [0:0] direct_interc_141_out;
wire [0:0] direct_interc_142_out;
wire [0:0] direct_interc_143_out;
wire [0:0] direct_interc_144_out;
wire [0:0] direct_interc_145_out;
wire [0:0] direct_interc_146_out;
wire [0:0] direct_interc_147_out;
wire [0:0] direct_interc_148_out;
wire [0:0] direct_interc_149_out;
wire [0:0] direct_interc_14_out;
wire [0:0] direct_interc_150_out;
wire [0:0] direct_interc_151_out;
wire [0:0] direct_interc_152_out;
wire [0:0] direct_interc_153_out;
wire [0:0] direct_interc_154_out;
wire [0:0] direct_interc_155_out;
wire [0:0] direct_interc_156_out;
wire [0:0] direct_interc_157_out;
wire [0:0] direct_interc_158_out;
wire [0:0] direct_interc_159_out;
wire [0:0] direct_interc_15_out;
wire [0:0] direct_interc_160_out;
wire [0:0] direct_interc_161_out;
wire [0:0] direct_interc_162_out;
wire [0:0] direct_interc_163_out;
wire [0:0] direct_interc_164_out;
wire [0:0] direct_interc_165_out;
wire [0:0] direct_interc_166_out;
wire [0:0] direct_interc_167_out;
wire [0:0] direct_interc_168_out;
wire [0:0] direct_interc_169_out;
wire [0:0] direct_interc_16_out;
wire [0:0] direct_interc_170_out;
wire [0:0] direct_interc_171_out;
wire [0:0] direct_interc_172_out;
wire [0:0] direct_interc_173_out;
wire [0:0] direct_interc_174_out;
wire [0:0] direct_interc_175_out;
wire [0:0] direct_interc_176_out;
wire [0:0] direct_interc_177_out;
wire [0:0] direct_interc_178_out;
wire [0:0] direct_interc_179_out;
wire [0:0] direct_interc_17_out;
wire [0:0] direct_interc_180_out;
wire [0:0] direct_interc_181_out;
wire [0:0] direct_interc_182_out;
wire [0:0] direct_interc_183_out;
wire [0:0] direct_interc_184_out;
wire [0:0] direct_interc_185_out;
wire [0:0] direct_interc_186_out;
wire [0:0] direct_interc_187_out;
wire [0:0] direct_interc_188_out;
wire [0:0] direct_interc_189_out;
wire [0:0] direct_interc_18_out;
wire [0:0] direct_interc_190_out;
wire [0:0] direct_interc_191_out;
wire [0:0] direct_interc_192_out;
wire [0:0] direct_interc_193_out;
wire [0:0] direct_interc_194_out;
wire [0:0] direct_interc_195_out;
wire [0:0] direct_interc_196_out;
wire [0:0] direct_interc_197_out;
wire [0:0] direct_interc_198_out;
wire [0:0] direct_interc_199_out;
wire [0:0] direct_interc_19_out;
wire [0:0] direct_interc_1_out;
wire [0:0] direct_interc_200_out;
wire [0:0] direct_interc_201_out;
wire [0:0] direct_interc_202_out;
wire [0:0] direct_interc_203_out;
wire [0:0] direct_interc_204_out;
wire [0:0] direct_interc_205_out;
wire [0:0] direct_interc_206_out;
wire [0:0] direct_interc_207_out;
wire [0:0] direct_interc_208_out;
wire [0:0] direct_interc_209_out;
wire [0:0] direct_interc_20_out;
wire [0:0] direct_interc_210_out;
wire [0:0] direct_interc_211_out;
wire [0:0] direct_interc_212_out;
wire [0:0] direct_interc_213_out;
wire [0:0] direct_interc_214_out;
wire [0:0] direct_interc_215_out;
wire [0:0] direct_interc_216_out;
wire [0:0] direct_interc_217_out;
wire [0:0] direct_interc_218_out;
wire [0:0] direct_interc_219_out;
wire [0:0] direct_interc_21_out;
wire [0:0] direct_interc_220_out;
wire [0:0] direct_interc_221_out;
wire [0:0] direct_interc_222_out;
wire [0:0] direct_interc_223_out;
wire [0:0] direct_interc_224_out;
wire [0:0] direct_interc_225_out;
wire [0:0] direct_interc_226_out;
wire [0:0] direct_interc_227_out;
wire [0:0] direct_interc_228_out;
wire [0:0] direct_interc_229_out;
wire [0:0] direct_interc_22_out;
wire [0:0] direct_interc_230_out;
wire [0:0] direct_interc_231_out;
wire [0:0] direct_interc_232_out;
wire [0:0] direct_interc_233_out;
wire [0:0] direct_interc_234_out;
wire [0:0] direct_interc_235_out;
wire [0:0] direct_interc_236_out;
wire [0:0] direct_interc_237_out;
wire [0:0] direct_interc_238_out;
wire [0:0] direct_interc_239_out;
wire [0:0] direct_interc_23_out;
wire [0:0] direct_interc_240_out;
wire [0:0] direct_interc_241_out;
wire [0:0] direct_interc_242_out;
wire [0:0] direct_interc_243_out;
wire [0:0] direct_interc_244_out;
wire [0:0] direct_interc_245_out;
wire [0:0] direct_interc_246_out;
wire [0:0] direct_interc_247_out;
wire [0:0] direct_interc_248_out;
wire [0:0] direct_interc_249_out;
wire [0:0] direct_interc_24_out;
wire [0:0] direct_interc_250_out;
wire [0:0] direct_interc_251_out;
wire [0:0] direct_interc_252_out;
wire [0:0] direct_interc_253_out;
wire [0:0] direct_interc_254_out;
wire [0:0] direct_interc_255_out;
wire [0:0] direct_interc_256_out;
wire [0:0] direct_interc_257_out;
wire [0:0] direct_interc_258_out;
wire [0:0] direct_interc_259_out;
wire [0:0] direct_interc_25_out;
wire [0:0] direct_interc_260_out;
wire [0:0] direct_interc_261_out;
wire [0:0] direct_interc_262_out;
wire [0:0] direct_interc_263_out;
wire [0:0] direct_interc_264_out;
wire [0:0] direct_interc_265_out;
wire [0:0] direct_interc_266_out;
wire [0:0] direct_interc_267_out;
wire [0:0] direct_interc_268_out;
wire [0:0] direct_interc_269_out;
wire [0:0] direct_interc_26_out;
wire [0:0] direct_interc_270_out;
wire [0:0] direct_interc_271_out;
wire [0:0] direct_interc_272_out;
wire [0:0] direct_interc_273_out;
wire [0:0] direct_interc_274_out;
wire [0:0] direct_interc_275_out;
wire [0:0] direct_interc_276_out;
wire [0:0] direct_interc_277_out;
wire [0:0] direct_interc_278_out;
wire [0:0] direct_interc_279_out;
wire [0:0] direct_interc_27_out;
wire [0:0] direct_interc_280_out;
wire [0:0] direct_interc_281_out;
wire [0:0] direct_interc_282_out;
wire [0:0] direct_interc_283_out;
wire [0:0] direct_interc_284_out;
wire [0:0] direct_interc_285_out;
wire [0:0] direct_interc_286_out;
wire [0:0] direct_interc_287_out;
wire [0:0] direct_interc_288_out;
wire [0:0] direct_interc_289_out;
wire [0:0] direct_interc_28_out;
wire [0:0] direct_interc_290_out;
wire [0:0] direct_interc_291_out;
wire [0:0] direct_interc_292_out;
wire [0:0] direct_interc_293_out;
wire [0:0] direct_interc_294_out;
wire [0:0] direct_interc_295_out;
wire [0:0] direct_interc_296_out;
wire [0:0] direct_interc_297_out;
wire [0:0] direct_interc_298_out;
wire [0:0] direct_interc_299_out;
wire [0:0] direct_interc_29_out;
wire [0:0] direct_interc_2_out;
wire [0:0] direct_interc_300_out;
wire [0:0] direct_interc_301_out;
wire [0:0] direct_interc_302_out;
wire [0:0] direct_interc_303_out;
wire [0:0] direct_interc_304_out;
wire [0:0] direct_interc_305_out;
wire [0:0] direct_interc_306_out;
wire [0:0] direct_interc_307_out;
wire [0:0] direct_interc_308_out;
wire [0:0] direct_interc_309_out;
wire [0:0] direct_interc_30_out;
wire [0:0] direct_interc_310_out;
wire [0:0] direct_interc_311_out;
wire [0:0] direct_interc_312_out;
wire [0:0] direct_interc_313_out;
wire [0:0] direct_interc_314_out;
wire [0:0] direct_interc_315_out;
wire [0:0] direct_interc_316_out;
wire [0:0] direct_interc_317_out;
wire [0:0] direct_interc_318_out;
wire [0:0] direct_interc_319_out;
wire [0:0] direct_interc_31_out;
wire [0:0] direct_interc_320_out;
wire [0:0] direct_interc_321_out;
wire [0:0] direct_interc_322_out;
wire [0:0] direct_interc_323_out;
wire [0:0] direct_interc_324_out;
wire [0:0] direct_interc_325_out;
wire [0:0] direct_interc_326_out;
wire [0:0] direct_interc_327_out;
wire [0:0] direct_interc_328_out;
wire [0:0] direct_interc_329_out;
wire [0:0] direct_interc_32_out;
wire [0:0] direct_interc_330_out;
wire [0:0] direct_interc_331_out;
wire [0:0] direct_interc_332_out;
wire [0:0] direct_interc_333_out;
wire [0:0] direct_interc_334_out;
wire [0:0] direct_interc_335_out;
wire [0:0] direct_interc_336_out;
wire [0:0] direct_interc_337_out;
wire [0:0] direct_interc_338_out;
wire [0:0] direct_interc_339_out;
wire [0:0] direct_interc_33_out;
wire [0:0] direct_interc_340_out;
wire [0:0] direct_interc_341_out;
wire [0:0] direct_interc_342_out;
wire [0:0] direct_interc_343_out;
wire [0:0] direct_interc_344_out;
wire [0:0] direct_interc_345_out;
wire [0:0] direct_interc_346_out;
wire [0:0] direct_interc_347_out;
wire [0:0] direct_interc_348_out;
wire [0:0] direct_interc_349_out;
wire [0:0] direct_interc_34_out;
wire [0:0] direct_interc_350_out;
wire [0:0] direct_interc_351_out;
wire [0:0] direct_interc_352_out;
wire [0:0] direct_interc_353_out;
wire [0:0] direct_interc_354_out;
wire [0:0] direct_interc_355_out;
wire [0:0] direct_interc_356_out;
wire [0:0] direct_interc_357_out;
wire [0:0] direct_interc_358_out;
wire [0:0] direct_interc_359_out;
wire [0:0] direct_interc_35_out;
wire [0:0] direct_interc_360_out;
wire [0:0] direct_interc_361_out;
wire [0:0] direct_interc_362_out;
wire [0:0] direct_interc_363_out;
wire [0:0] direct_interc_364_out;
wire [0:0] direct_interc_365_out;
wire [0:0] direct_interc_366_out;
wire [0:0] direct_interc_367_out;
wire [0:0] direct_interc_368_out;
wire [0:0] direct_interc_369_out;
wire [0:0] direct_interc_36_out;
wire [0:0] direct_interc_370_out;
wire [0:0] direct_interc_371_out;
wire [0:0] direct_interc_372_out;
wire [0:0] direct_interc_373_out;
wire [0:0] direct_interc_374_out;
wire [0:0] direct_interc_375_out;
wire [0:0] direct_interc_376_out;
wire [0:0] direct_interc_377_out;
wire [0:0] direct_interc_378_out;
wire [0:0] direct_interc_379_out;
wire [0:0] direct_interc_37_out;
wire [0:0] direct_interc_380_out;
wire [0:0] direct_interc_381_out;
wire [0:0] direct_interc_382_out;
wire [0:0] direct_interc_383_out;
wire [0:0] direct_interc_384_out;
wire [0:0] direct_interc_385_out;
wire [0:0] direct_interc_386_out;
wire [0:0] direct_interc_387_out;
wire [0:0] direct_interc_388_out;
wire [0:0] direct_interc_389_out;
wire [0:0] direct_interc_38_out;
wire [0:0] direct_interc_390_out;
wire [0:0] direct_interc_391_out;
wire [0:0] direct_interc_392_out;
wire [0:0] direct_interc_393_out;
wire [0:0] direct_interc_394_out;
wire [0:0] direct_interc_395_out;
wire [0:0] direct_interc_396_out;
wire [0:0] direct_interc_397_out;
wire [0:0] direct_interc_398_out;
wire [0:0] direct_interc_399_out;
wire [0:0] direct_interc_39_out;
wire [0:0] direct_interc_3_out;
wire [0:0] direct_interc_400_out;
wire [0:0] direct_interc_401_out;
wire [0:0] direct_interc_402_out;
wire [0:0] direct_interc_403_out;
wire [0:0] direct_interc_404_out;
wire [0:0] direct_interc_405_out;
wire [0:0] direct_interc_406_out;
wire [0:0] direct_interc_407_out;
wire [0:0] direct_interc_408_out;
wire [0:0] direct_interc_409_out;
wire [0:0] direct_interc_40_out;
wire [0:0] direct_interc_410_out;
wire [0:0] direct_interc_411_out;
wire [0:0] direct_interc_412_out;
wire [0:0] direct_interc_413_out;
wire [0:0] direct_interc_414_out;
wire [0:0] direct_interc_415_out;
wire [0:0] direct_interc_416_out;
wire [0:0] direct_interc_417_out;
wire [0:0] direct_interc_418_out;
wire [0:0] direct_interc_419_out;
wire [0:0] direct_interc_41_out;
wire [0:0] direct_interc_420_out;
wire [0:0] direct_interc_421_out;
wire [0:0] direct_interc_422_out;
wire [0:0] direct_interc_423_out;
wire [0:0] direct_interc_424_out;
wire [0:0] direct_interc_425_out;
wire [0:0] direct_interc_426_out;
wire [0:0] direct_interc_427_out;
wire [0:0] direct_interc_428_out;
wire [0:0] direct_interc_429_out;
wire [0:0] direct_interc_42_out;
wire [0:0] direct_interc_430_out;
wire [0:0] direct_interc_431_out;
wire [0:0] direct_interc_432_out;
wire [0:0] direct_interc_433_out;
wire [0:0] direct_interc_434_out;
wire [0:0] direct_interc_435_out;
wire [0:0] direct_interc_436_out;
wire [0:0] direct_interc_437_out;
wire [0:0] direct_interc_438_out;
wire [0:0] direct_interc_439_out;
wire [0:0] direct_interc_43_out;
wire [0:0] direct_interc_440_out;
wire [0:0] direct_interc_441_out;
wire [0:0] direct_interc_442_out;
wire [0:0] direct_interc_443_out;
wire [0:0] direct_interc_444_out;
wire [0:0] direct_interc_445_out;
wire [0:0] direct_interc_446_out;
wire [0:0] direct_interc_447_out;
wire [0:0] direct_interc_448_out;
wire [0:0] direct_interc_449_out;
wire [0:0] direct_interc_44_out;
wire [0:0] direct_interc_450_out;
wire [0:0] direct_interc_451_out;
wire [0:0] direct_interc_452_out;
wire [0:0] direct_interc_453_out;
wire [0:0] direct_interc_454_out;
wire [0:0] direct_interc_455_out;
wire [0:0] direct_interc_456_out;
wire [0:0] direct_interc_457_out;
wire [0:0] direct_interc_458_out;
wire [0:0] direct_interc_459_out;
wire [0:0] direct_interc_45_out;
wire [0:0] direct_interc_460_out;
wire [0:0] direct_interc_461_out;
wire [0:0] direct_interc_462_out;
wire [0:0] direct_interc_463_out;
wire [0:0] direct_interc_464_out;
wire [0:0] direct_interc_465_out;
wire [0:0] direct_interc_466_out;
wire [0:0] direct_interc_467_out;
wire [0:0] direct_interc_468_out;
wire [0:0] direct_interc_469_out;
wire [0:0] direct_interc_46_out;
wire [0:0] direct_interc_470_out;
wire [0:0] direct_interc_471_out;
wire [0:0] direct_interc_472_out;
wire [0:0] direct_interc_473_out;
wire [0:0] direct_interc_474_out;
wire [0:0] direct_interc_475_out;
wire [0:0] direct_interc_476_out;
wire [0:0] direct_interc_477_out;
wire [0:0] direct_interc_478_out;
wire [0:0] direct_interc_479_out;
wire [0:0] direct_interc_47_out;
wire [0:0] direct_interc_480_out;
wire [0:0] direct_interc_481_out;
wire [0:0] direct_interc_482_out;
wire [0:0] direct_interc_483_out;
wire [0:0] direct_interc_484_out;
wire [0:0] direct_interc_485_out;
wire [0:0] direct_interc_486_out;
wire [0:0] direct_interc_487_out;
wire [0:0] direct_interc_488_out;
wire [0:0] direct_interc_489_out;
wire [0:0] direct_interc_48_out;
wire [0:0] direct_interc_490_out;
wire [0:0] direct_interc_491_out;
wire [0:0] direct_interc_492_out;
wire [0:0] direct_interc_493_out;
wire [0:0] direct_interc_494_out;
wire [0:0] direct_interc_495_out;
wire [0:0] direct_interc_496_out;
wire [0:0] direct_interc_497_out;
wire [0:0] direct_interc_498_out;
wire [0:0] direct_interc_499_out;
wire [0:0] direct_interc_49_out;
wire [0:0] direct_interc_4_out;
wire [0:0] direct_interc_500_out;
wire [0:0] direct_interc_501_out;
wire [0:0] direct_interc_502_out;
wire [0:0] direct_interc_503_out;
wire [0:0] direct_interc_504_out;
wire [0:0] direct_interc_505_out;
wire [0:0] direct_interc_506_out;
wire [0:0] direct_interc_507_out;
wire [0:0] direct_interc_508_out;
wire [0:0] direct_interc_509_out;
wire [0:0] direct_interc_50_out;
wire [0:0] direct_interc_510_out;
wire [0:0] direct_interc_511_out;
wire [0:0] direct_interc_512_out;
wire [0:0] direct_interc_513_out;
wire [0:0] direct_interc_514_out;
wire [0:0] direct_interc_515_out;
wire [0:0] direct_interc_516_out;
wire [0:0] direct_interc_517_out;
wire [0:0] direct_interc_518_out;
wire [0:0] direct_interc_519_out;
wire [0:0] direct_interc_51_out;
wire [0:0] direct_interc_520_out;
wire [0:0] direct_interc_521_out;
wire [0:0] direct_interc_522_out;
wire [0:0] direct_interc_523_out;
wire [0:0] direct_interc_524_out;
wire [0:0] direct_interc_525_out;
wire [0:0] direct_interc_526_out;
wire [0:0] direct_interc_527_out;
wire [0:0] direct_interc_528_out;
wire [0:0] direct_interc_529_out;
wire [0:0] direct_interc_52_out;
wire [0:0] direct_interc_530_out;
wire [0:0] direct_interc_531_out;
wire [0:0] direct_interc_532_out;
wire [0:0] direct_interc_533_out;
wire [0:0] direct_interc_534_out;
wire [0:0] direct_interc_535_out;
wire [0:0] direct_interc_536_out;
wire [0:0] direct_interc_537_out;
wire [0:0] direct_interc_538_out;
wire [0:0] direct_interc_539_out;
wire [0:0] direct_interc_53_out;
wire [0:0] direct_interc_540_out;
wire [0:0] direct_interc_541_out;
wire [0:0] direct_interc_542_out;
wire [0:0] direct_interc_543_out;
wire [0:0] direct_interc_544_out;
wire [0:0] direct_interc_545_out;
wire [0:0] direct_interc_546_out;
wire [0:0] direct_interc_547_out;
wire [0:0] direct_interc_548_out;
wire [0:0] direct_interc_549_out;
wire [0:0] direct_interc_54_out;
wire [0:0] direct_interc_550_out;
wire [0:0] direct_interc_551_out;
wire [0:0] direct_interc_552_out;
wire [0:0] direct_interc_553_out;
wire [0:0] direct_interc_554_out;
wire [0:0] direct_interc_555_out;
wire [0:0] direct_interc_556_out;
wire [0:0] direct_interc_557_out;
wire [0:0] direct_interc_558_out;
wire [0:0] direct_interc_559_out;
wire [0:0] direct_interc_55_out;
wire [0:0] direct_interc_560_out;
wire [0:0] direct_interc_561_out;
wire [0:0] direct_interc_562_out;
wire [0:0] direct_interc_563_out;
wire [0:0] direct_interc_564_out;
wire [0:0] direct_interc_565_out;
wire [0:0] direct_interc_566_out;
wire [0:0] direct_interc_567_out;
wire [0:0] direct_interc_568_out;
wire [0:0] direct_interc_569_out;
wire [0:0] direct_interc_56_out;
wire [0:0] direct_interc_570_out;
wire [0:0] direct_interc_571_out;
wire [0:0] direct_interc_572_out;
wire [0:0] direct_interc_573_out;
wire [0:0] direct_interc_574_out;
wire [0:0] direct_interc_575_out;
wire [0:0] direct_interc_576_out;
wire [0:0] direct_interc_577_out;
wire [0:0] direct_interc_578_out;
wire [0:0] direct_interc_579_out;
wire [0:0] direct_interc_57_out;
wire [0:0] direct_interc_580_out;
wire [0:0] direct_interc_581_out;
wire [0:0] direct_interc_582_out;
wire [0:0] direct_interc_583_out;
wire [0:0] direct_interc_584_out;
wire [0:0] direct_interc_585_out;
wire [0:0] direct_interc_586_out;
wire [0:0] direct_interc_587_out;
wire [0:0] direct_interc_588_out;
wire [0:0] direct_interc_589_out;
wire [0:0] direct_interc_58_out;
wire [0:0] direct_interc_590_out;
wire [0:0] direct_interc_591_out;
wire [0:0] direct_interc_592_out;
wire [0:0] direct_interc_593_out;
wire [0:0] direct_interc_594_out;
wire [0:0] direct_interc_595_out;
wire [0:0] direct_interc_596_out;
wire [0:0] direct_interc_597_out;
wire [0:0] direct_interc_598_out;
wire [0:0] direct_interc_599_out;
wire [0:0] direct_interc_59_out;
wire [0:0] direct_interc_5_out;
wire [0:0] direct_interc_600_out;
wire [0:0] direct_interc_601_out;
wire [0:0] direct_interc_602_out;
wire [0:0] direct_interc_603_out;
wire [0:0] direct_interc_604_out;
wire [0:0] direct_interc_605_out;
wire [0:0] direct_interc_606_out;
wire [0:0] direct_interc_607_out;
wire [0:0] direct_interc_608_out;
wire [0:0] direct_interc_609_out;
wire [0:0] direct_interc_60_out;
wire [0:0] direct_interc_610_out;
wire [0:0] direct_interc_611_out;
wire [0:0] direct_interc_612_out;
wire [0:0] direct_interc_613_out;
wire [0:0] direct_interc_614_out;
wire [0:0] direct_interc_615_out;
wire [0:0] direct_interc_616_out;
wire [0:0] direct_interc_617_out;
wire [0:0] direct_interc_618_out;
wire [0:0] direct_interc_619_out;
wire [0:0] direct_interc_61_out;
wire [0:0] direct_interc_620_out;
wire [0:0] direct_interc_621_out;
wire [0:0] direct_interc_622_out;
wire [0:0] direct_interc_623_out;
wire [0:0] direct_interc_624_out;
wire [0:0] direct_interc_625_out;
wire [0:0] direct_interc_626_out;
wire [0:0] direct_interc_627_out;
wire [0:0] direct_interc_628_out;
wire [0:0] direct_interc_629_out;
wire [0:0] direct_interc_62_out;
wire [0:0] direct_interc_630_out;
wire [0:0] direct_interc_631_out;
wire [0:0] direct_interc_632_out;
wire [0:0] direct_interc_633_out;
wire [0:0] direct_interc_634_out;
wire [0:0] direct_interc_635_out;
wire [0:0] direct_interc_636_out;
wire [0:0] direct_interc_637_out;
wire [0:0] direct_interc_638_out;
wire [0:0] direct_interc_639_out;
wire [0:0] direct_interc_63_out;
wire [0:0] direct_interc_640_out;
wire [0:0] direct_interc_641_out;
wire [0:0] direct_interc_642_out;
wire [0:0] direct_interc_643_out;
wire [0:0] direct_interc_644_out;
wire [0:0] direct_interc_645_out;
wire [0:0] direct_interc_646_out;
wire [0:0] direct_interc_647_out;
wire [0:0] direct_interc_648_out;
wire [0:0] direct_interc_649_out;
wire [0:0] direct_interc_64_out;
wire [0:0] direct_interc_650_out;
wire [0:0] direct_interc_651_out;
wire [0:0] direct_interc_652_out;
wire [0:0] direct_interc_653_out;
wire [0:0] direct_interc_654_out;
wire [0:0] direct_interc_655_out;
wire [0:0] direct_interc_656_out;
wire [0:0] direct_interc_657_out;
wire [0:0] direct_interc_658_out;
wire [0:0] direct_interc_659_out;
wire [0:0] direct_interc_65_out;
wire [0:0] direct_interc_660_out;
wire [0:0] direct_interc_661_out;
wire [0:0] direct_interc_662_out;
wire [0:0] direct_interc_663_out;
wire [0:0] direct_interc_664_out;
wire [0:0] direct_interc_665_out;
wire [0:0] direct_interc_666_out;
wire [0:0] direct_interc_667_out;
wire [0:0] direct_interc_668_out;
wire [0:0] direct_interc_669_out;
wire [0:0] direct_interc_66_out;
wire [0:0] direct_interc_670_out;
wire [0:0] direct_interc_671_out;
wire [0:0] direct_interc_672_out;
wire [0:0] direct_interc_673_out;
wire [0:0] direct_interc_674_out;
wire [0:0] direct_interc_675_out;
wire [0:0] direct_interc_676_out;
wire [0:0] direct_interc_677_out;
wire [0:0] direct_interc_678_out;
wire [0:0] direct_interc_679_out;
wire [0:0] direct_interc_67_out;
wire [0:0] direct_interc_680_out;
wire [0:0] direct_interc_681_out;
wire [0:0] direct_interc_682_out;
wire [0:0] direct_interc_683_out;
wire [0:0] direct_interc_684_out;
wire [0:0] direct_interc_685_out;
wire [0:0] direct_interc_686_out;
wire [0:0] direct_interc_687_out;
wire [0:0] direct_interc_688_out;
wire [0:0] direct_interc_689_out;
wire [0:0] direct_interc_68_out;
wire [0:0] direct_interc_690_out;
wire [0:0] direct_interc_691_out;
wire [0:0] direct_interc_692_out;
wire [0:0] direct_interc_693_out;
wire [0:0] direct_interc_694_out;
wire [0:0] direct_interc_695_out;
wire [0:0] direct_interc_696_out;
wire [0:0] direct_interc_697_out;
wire [0:0] direct_interc_698_out;
wire [0:0] direct_interc_699_out;
wire [0:0] direct_interc_69_out;
wire [0:0] direct_interc_6_out;
wire [0:0] direct_interc_700_out;
wire [0:0] direct_interc_701_out;
wire [0:0] direct_interc_702_out;
wire [0:0] direct_interc_703_out;
wire [0:0] direct_interc_704_out;
wire [0:0] direct_interc_705_out;
wire [0:0] direct_interc_706_out;
wire [0:0] direct_interc_707_out;
wire [0:0] direct_interc_708_out;
wire [0:0] direct_interc_709_out;
wire [0:0] direct_interc_70_out;
wire [0:0] direct_interc_710_out;
wire [0:0] direct_interc_711_out;
wire [0:0] direct_interc_712_out;
wire [0:0] direct_interc_713_out;
wire [0:0] direct_interc_714_out;
wire [0:0] direct_interc_715_out;
wire [0:0] direct_interc_716_out;
wire [0:0] direct_interc_717_out;
wire [0:0] direct_interc_718_out;
wire [0:0] direct_interc_719_out;
wire [0:0] direct_interc_71_out;
wire [0:0] direct_interc_720_out;
wire [0:0] direct_interc_721_out;
wire [0:0] direct_interc_722_out;
wire [0:0] direct_interc_723_out;
wire [0:0] direct_interc_724_out;
wire [0:0] direct_interc_725_out;
wire [0:0] direct_interc_726_out;
wire [0:0] direct_interc_727_out;
wire [0:0] direct_interc_728_out;
wire [0:0] direct_interc_729_out;
wire [0:0] direct_interc_72_out;
wire [0:0] direct_interc_730_out;
wire [0:0] direct_interc_731_out;
wire [0:0] direct_interc_732_out;
wire [0:0] direct_interc_733_out;
wire [0:0] direct_interc_734_out;
wire [0:0] direct_interc_735_out;
wire [0:0] direct_interc_736_out;
wire [0:0] direct_interc_737_out;
wire [0:0] direct_interc_738_out;
wire [0:0] direct_interc_739_out;
wire [0:0] direct_interc_73_out;
wire [0:0] direct_interc_740_out;
wire [0:0] direct_interc_741_out;
wire [0:0] direct_interc_742_out;
wire [0:0] direct_interc_743_out;
wire [0:0] direct_interc_744_out;
wire [0:0] direct_interc_745_out;
wire [0:0] direct_interc_746_out;
wire [0:0] direct_interc_747_out;
wire [0:0] direct_interc_748_out;
wire [0:0] direct_interc_749_out;
wire [0:0] direct_interc_74_out;
wire [0:0] direct_interc_750_out;
wire [0:0] direct_interc_751_out;
wire [0:0] direct_interc_752_out;
wire [0:0] direct_interc_753_out;
wire [0:0] direct_interc_754_out;
wire [0:0] direct_interc_755_out;
wire [0:0] direct_interc_756_out;
wire [0:0] direct_interc_757_out;
wire [0:0] direct_interc_758_out;
wire [0:0] direct_interc_759_out;
wire [0:0] direct_interc_75_out;
wire [0:0] direct_interc_760_out;
wire [0:0] direct_interc_761_out;
wire [0:0] direct_interc_762_out;
wire [0:0] direct_interc_763_out;
wire [0:0] direct_interc_764_out;
wire [0:0] direct_interc_765_out;
wire [0:0] direct_interc_766_out;
wire [0:0] direct_interc_767_out;
wire [0:0] direct_interc_768_out;
wire [0:0] direct_interc_769_out;
wire [0:0] direct_interc_76_out;
wire [0:0] direct_interc_770_out;
wire [0:0] direct_interc_771_out;
wire [0:0] direct_interc_772_out;
wire [0:0] direct_interc_773_out;
wire [0:0] direct_interc_774_out;
wire [0:0] direct_interc_775_out;
wire [0:0] direct_interc_776_out;
wire [0:0] direct_interc_777_out;
wire [0:0] direct_interc_778_out;
wire [0:0] direct_interc_779_out;
wire [0:0] direct_interc_77_out;
wire [0:0] direct_interc_780_out;
wire [0:0] direct_interc_781_out;
wire [0:0] direct_interc_782_out;
wire [0:0] direct_interc_783_out;
wire [0:0] direct_interc_784_out;
wire [0:0] direct_interc_785_out;
wire [0:0] direct_interc_786_out;
wire [0:0] direct_interc_787_out;
wire [0:0] direct_interc_788_out;
wire [0:0] direct_interc_789_out;
wire [0:0] direct_interc_78_out;
wire [0:0] direct_interc_790_out;
wire [0:0] direct_interc_791_out;
wire [0:0] direct_interc_792_out;
wire [0:0] direct_interc_793_out;
wire [0:0] direct_interc_794_out;
wire [0:0] direct_interc_795_out;
wire [0:0] direct_interc_796_out;
wire [0:0] direct_interc_797_out;
wire [0:0] direct_interc_798_out;
wire [0:0] direct_interc_799_out;
wire [0:0] direct_interc_79_out;
wire [0:0] direct_interc_7_out;
wire [0:0] direct_interc_800_out;
wire [0:0] direct_interc_801_out;
wire [0:0] direct_interc_802_out;
wire [0:0] direct_interc_803_out;
wire [0:0] direct_interc_804_out;
wire [0:0] direct_interc_805_out;
wire [0:0] direct_interc_806_out;
wire [0:0] direct_interc_807_out;
wire [0:0] direct_interc_808_out;
wire [0:0] direct_interc_809_out;
wire [0:0] direct_interc_80_out;
wire [0:0] direct_interc_810_out;
wire [0:0] direct_interc_811_out;
wire [0:0] direct_interc_812_out;
wire [0:0] direct_interc_813_out;
wire [0:0] direct_interc_814_out;
wire [0:0] direct_interc_815_out;
wire [0:0] direct_interc_816_out;
wire [0:0] direct_interc_817_out;
wire [0:0] direct_interc_818_out;
wire [0:0] direct_interc_819_out;
wire [0:0] direct_interc_81_out;
wire [0:0] direct_interc_820_out;
wire [0:0] direct_interc_821_out;
wire [0:0] direct_interc_822_out;
wire [0:0] direct_interc_823_out;
wire [0:0] direct_interc_824_out;
wire [0:0] direct_interc_825_out;
wire [0:0] direct_interc_826_out;
wire [0:0] direct_interc_827_out;
wire [0:0] direct_interc_828_out;
wire [0:0] direct_interc_829_out;
wire [0:0] direct_interc_82_out;
wire [0:0] direct_interc_830_out;
wire [0:0] direct_interc_831_out;
wire [0:0] direct_interc_832_out;
wire [0:0] direct_interc_833_out;
wire [0:0] direct_interc_834_out;
wire [0:0] direct_interc_835_out;
wire [0:0] direct_interc_836_out;
wire [0:0] direct_interc_837_out;
wire [0:0] direct_interc_838_out;
wire [0:0] direct_interc_839_out;
wire [0:0] direct_interc_83_out;
wire [0:0] direct_interc_840_out;
wire [0:0] direct_interc_841_out;
wire [0:0] direct_interc_842_out;
wire [0:0] direct_interc_843_out;
wire [0:0] direct_interc_844_out;
wire [0:0] direct_interc_845_out;
wire [0:0] direct_interc_846_out;
wire [0:0] direct_interc_847_out;
wire [0:0] direct_interc_848_out;
wire [0:0] direct_interc_849_out;
wire [0:0] direct_interc_84_out;
wire [0:0] direct_interc_85_out;
wire [0:0] direct_interc_86_out;
wire [0:0] direct_interc_87_out;
wire [0:0] direct_interc_88_out;
wire [0:0] direct_interc_89_out;
wire [0:0] direct_interc_8_out;
wire [0:0] direct_interc_90_out;
wire [0:0] direct_interc_91_out;
wire [0:0] direct_interc_92_out;
wire [0:0] direct_interc_93_out;
wire [0:0] direct_interc_94_out;
wire [0:0] direct_interc_95_out;
wire [0:0] direct_interc_96_out;
wire [0:0] direct_interc_97_out;
wire [0:0] direct_interc_98_out;
wire [0:0] direct_interc_99_out;
wire [0:0] direct_interc_9_out;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_0_ff_IACK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_1_ff_IACK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_0_ff_IACK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_1_ff_IACK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_0_ff_IACK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_1_ff_IACK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_0_ff_IACK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_1_ff_IACK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_0_ff_IACK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_1_ff_IACK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_0_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_10_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_11_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_12_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_13_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_14_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_15_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_16_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_17_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_18_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_19_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_1_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_20_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_21_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_22_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_23_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_24_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_25_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_26_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_27_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_28_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_29_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_2_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_30_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_31_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_32_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_33_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_34_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_3_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_4_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_5_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_6_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_7_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_8_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_9_ff_IDATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_0_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_10_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_11_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_12_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_13_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_14_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_15_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_16_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_17_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_18_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_19_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_1_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_20_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_21_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_22_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_23_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_24_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_25_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_26_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_27_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_28_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_29_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_2_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_30_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_31_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_32_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_33_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_34_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_3_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_4_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_5_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_6_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_7_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_8_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_9_ff_IDATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_0_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_10_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_11_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_12_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_13_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_14_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_15_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_16_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_17_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_18_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_19_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_1_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_20_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_21_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_22_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_23_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_24_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_25_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_26_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_27_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_28_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_29_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_2_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_30_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_31_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_32_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_33_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_34_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_3_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_4_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_5_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_6_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_7_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_8_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_9_ff_IDATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_0_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_10_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_11_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_12_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_13_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_14_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_15_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_16_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_17_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_18_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_19_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_1_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_20_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_21_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_22_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_23_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_24_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_25_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_26_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_27_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_28_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_29_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_2_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_30_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_31_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_32_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_33_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_34_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_3_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_4_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_5_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_6_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_7_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_8_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_9_ff_IDATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_0_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_10_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_11_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_12_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_13_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_14_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_15_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_16_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_17_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_18_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_19_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_1_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_20_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_21_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_22_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_23_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_24_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_25_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_26_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_27_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_28_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_29_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_2_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_30_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_31_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_32_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_33_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_34_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_3_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_4_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_5_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_6_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_7_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_8_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_9_ff_IDATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_0_ff_ILCK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_1_ff_ILCK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_0_ff_ILCK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_1_ff_ILCK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_0_ff_ILCK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_1_ff_ILCK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_0_ff_ILCK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_1_ff_ILCK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_0_ff_ILCK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_1_ff_ILCK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_0_0_ff_IVALID_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_1_0_ff_IVALID_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_2_0_ff_IVALID_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_3_0_ff_IVALID_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_4_0_ff_IVALID_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_0_0_ff_IVCH_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_1_0_ff_IVCH_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_2_0_ff_IVCH_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_3_0_ff_IVCH_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_4_0_ff_IVCH_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_0_ff_MY_XPOS_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_1_ff_MY_XPOS_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_0_ff_MY_YPOS_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_1_ff_MY_YPOS_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_0_ff_OACK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_1_ff_OACK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_0_ff_OACK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_1_ff_OACK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_0_ff_OACK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_1_ff_OACK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_0_ff_OACK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_1_ff_OACK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_0_ff_OACK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_1_ff_OACK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_0_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_10_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_11_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_12_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_13_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_14_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_15_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_16_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_17_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_18_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_19_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_1_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_20_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_21_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_22_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_23_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_24_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_25_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_26_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_27_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_28_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_29_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_2_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_30_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_31_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_32_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_33_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_34_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_3_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_4_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_5_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_6_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_7_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_8_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_9_ff_ODATA_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_0_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_10_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_11_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_12_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_13_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_14_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_15_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_16_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_17_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_18_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_19_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_1_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_20_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_21_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_22_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_23_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_24_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_25_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_26_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_27_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_28_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_29_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_2_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_30_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_31_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_32_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_33_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_34_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_3_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_4_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_5_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_6_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_7_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_8_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_9_ff_ODATA_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_0_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_10_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_11_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_12_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_13_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_14_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_15_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_16_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_17_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_18_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_19_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_1_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_20_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_21_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_22_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_23_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_24_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_25_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_26_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_27_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_28_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_29_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_2_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_30_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_31_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_32_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_33_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_34_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_3_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_4_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_5_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_6_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_7_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_8_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_9_ff_ODATA_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_0_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_10_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_11_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_12_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_13_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_14_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_15_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_16_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_17_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_18_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_19_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_1_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_20_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_21_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_22_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_23_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_24_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_25_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_26_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_27_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_28_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_29_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_2_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_30_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_31_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_32_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_33_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_34_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_3_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_4_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_5_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_6_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_7_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_8_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_9_ff_ODATA_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_0_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_10_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_11_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_12_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_13_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_14_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_15_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_16_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_17_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_18_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_19_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_1_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_20_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_21_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_22_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_23_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_24_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_25_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_26_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_27_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_28_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_29_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_2_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_30_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_31_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_32_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_33_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_34_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_3_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_4_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_5_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_6_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_7_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_8_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_9_ff_ODATA_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_0_ff_OLCK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_1_ff_OLCK_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_0_ff_OLCK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_1_ff_OLCK_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_0_ff_OLCK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_1_ff_OLCK_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_0_ff_OLCK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_1_ff_OLCK_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_0_ff_OLCK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_1_ff_OLCK_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_0_ff_ORDY_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_1_ff_ORDY_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_0_ff_ORDY_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_1_ff_ORDY_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_0_ff_ORDY_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_1_ff_ORDY_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_0_ff_ORDY_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_1_ff_ORDY_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_0_ff_ORDY_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_1_ff_ORDY_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_0_0_ff_OVALID_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_1_0_ff_OVALID_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_2_0_ff_OVALID_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_3_0_ff_OVALID_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_4_0_ff_OVALID_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_0_0_ff_OVCH_0_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_1_0_ff_OVCH_1_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_2_0_ff_OVCH_2_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_3_0_ff_OVCH_3_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_4_0_ff_OVCH_4_Q;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_RST__0_ff_RST__Q;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4;
wire [0:34] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0;
wire [0:34] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1;
wire [0:34] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2;
wire [0:34] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3;
wire [0:34] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3;
wire [0:1] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_0;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_1;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_2;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_3;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_4;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_0;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_1;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_2;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_3;
wire [0:0] logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_4;
wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_100_sram;
wire [0:1] mux_tree_tapbuf_size2_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_101_sram;
wire [0:1] mux_tree_tapbuf_size2_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_102_sram;
wire [0:1] mux_tree_tapbuf_size2_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_103_sram;
wire [0:1] mux_tree_tapbuf_size2_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_104_sram;
wire [0:1] mux_tree_tapbuf_size2_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_105_sram;
wire [0:1] mux_tree_tapbuf_size2_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_106_sram;
wire [0:1] mux_tree_tapbuf_size2_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_107_sram;
wire [0:1] mux_tree_tapbuf_size2_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_108_sram;
wire [0:1] mux_tree_tapbuf_size2_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_109_sram;
wire [0:1] mux_tree_tapbuf_size2_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_110_sram;
wire [0:1] mux_tree_tapbuf_size2_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_111_sram;
wire [0:1] mux_tree_tapbuf_size2_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_112_sram;
wire [0:1] mux_tree_tapbuf_size2_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_113_sram;
wire [0:1] mux_tree_tapbuf_size2_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_114_sram;
wire [0:1] mux_tree_tapbuf_size2_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_115_sram;
wire [0:1] mux_tree_tapbuf_size2_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_116_sram;
wire [0:1] mux_tree_tapbuf_size2_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_117_sram;
wire [0:1] mux_tree_tapbuf_size2_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_118_sram;
wire [0:1] mux_tree_tapbuf_size2_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_119_sram;
wire [0:1] mux_tree_tapbuf_size2_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_120_sram;
wire [0:1] mux_tree_tapbuf_size2_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_121_sram;
wire [0:1] mux_tree_tapbuf_size2_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_122_sram;
wire [0:1] mux_tree_tapbuf_size2_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_123_sram;
wire [0:1] mux_tree_tapbuf_size2_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_124_sram;
wire [0:1] mux_tree_tapbuf_size2_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_125_sram;
wire [0:1] mux_tree_tapbuf_size2_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_126_sram;
wire [0:1] mux_tree_tapbuf_size2_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_127_sram;
wire [0:1] mux_tree_tapbuf_size2_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_128_sram;
wire [0:1] mux_tree_tapbuf_size2_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_129_sram;
wire [0:1] mux_tree_tapbuf_size2_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_130_sram;
wire [0:1] mux_tree_tapbuf_size2_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_131_sram;
wire [0:1] mux_tree_tapbuf_size2_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_132_sram;
wire [0:1] mux_tree_tapbuf_size2_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_133_sram;
wire [0:1] mux_tree_tapbuf_size2_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_134_sram;
wire [0:1] mux_tree_tapbuf_size2_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_135_sram;
wire [0:1] mux_tree_tapbuf_size2_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_136_sram;
wire [0:1] mux_tree_tapbuf_size2_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_137_sram;
wire [0:1] mux_tree_tapbuf_size2_137_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_138_sram;
wire [0:1] mux_tree_tapbuf_size2_138_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_139_sram;
wire [0:1] mux_tree_tapbuf_size2_139_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_140_sram;
wire [0:1] mux_tree_tapbuf_size2_140_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_141_sram;
wire [0:1] mux_tree_tapbuf_size2_141_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_142_sram;
wire [0:1] mux_tree_tapbuf_size2_142_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_143_sram;
wire [0:1] mux_tree_tapbuf_size2_143_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_144_sram;
wire [0:1] mux_tree_tapbuf_size2_144_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_145_sram;
wire [0:1] mux_tree_tapbuf_size2_145_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_146_sram;
wire [0:1] mux_tree_tapbuf_size2_146_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_147_sram;
wire [0:1] mux_tree_tapbuf_size2_147_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_148_sram;
wire [0:1] mux_tree_tapbuf_size2_148_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_149_sram;
wire [0:1] mux_tree_tapbuf_size2_149_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_150_sram;
wire [0:1] mux_tree_tapbuf_size2_150_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_151_sram;
wire [0:1] mux_tree_tapbuf_size2_151_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_152_sram;
wire [0:1] mux_tree_tapbuf_size2_152_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_153_sram;
wire [0:1] mux_tree_tapbuf_size2_153_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_154_sram;
wire [0:1] mux_tree_tapbuf_size2_154_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_155_sram;
wire [0:1] mux_tree_tapbuf_size2_155_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_156_sram;
wire [0:1] mux_tree_tapbuf_size2_156_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_157_sram;
wire [0:1] mux_tree_tapbuf_size2_157_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_158_sram;
wire [0:1] mux_tree_tapbuf_size2_158_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_159_sram;
wire [0:1] mux_tree_tapbuf_size2_159_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_160_sram;
wire [0:1] mux_tree_tapbuf_size2_160_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_161_sram;
wire [0:1] mux_tree_tapbuf_size2_161_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_162_sram;
wire [0:1] mux_tree_tapbuf_size2_162_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_163_sram;
wire [0:1] mux_tree_tapbuf_size2_163_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_164_sram;
wire [0:1] mux_tree_tapbuf_size2_164_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_165_sram;
wire [0:1] mux_tree_tapbuf_size2_165_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_166_sram;
wire [0:1] mux_tree_tapbuf_size2_166_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_167_sram;
wire [0:1] mux_tree_tapbuf_size2_167_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_168_sram;
wire [0:1] mux_tree_tapbuf_size2_168_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_169_sram;
wire [0:1] mux_tree_tapbuf_size2_169_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_170_sram;
wire [0:1] mux_tree_tapbuf_size2_170_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_171_sram;
wire [0:1] mux_tree_tapbuf_size2_171_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_172_sram;
wire [0:1] mux_tree_tapbuf_size2_172_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_173_sram;
wire [0:1] mux_tree_tapbuf_size2_173_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_174_sram;
wire [0:1] mux_tree_tapbuf_size2_174_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_175_sram;
wire [0:1] mux_tree_tapbuf_size2_175_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_176_sram;
wire [0:1] mux_tree_tapbuf_size2_176_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_177_sram;
wire [0:1] mux_tree_tapbuf_size2_177_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_178_sram;
wire [0:1] mux_tree_tapbuf_size2_178_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_179_sram;
wire [0:1] mux_tree_tapbuf_size2_179_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_180_sram;
wire [0:1] mux_tree_tapbuf_size2_180_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_181_sram;
wire [0:1] mux_tree_tapbuf_size2_181_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_182_sram;
wire [0:1] mux_tree_tapbuf_size2_182_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_183_sram;
wire [0:1] mux_tree_tapbuf_size2_183_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_184_sram;
wire [0:1] mux_tree_tapbuf_size2_184_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_185_sram;
wire [0:1] mux_tree_tapbuf_size2_185_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_186_sram;
wire [0:1] mux_tree_tapbuf_size2_186_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_187_sram;
wire [0:1] mux_tree_tapbuf_size2_187_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_188_sram;
wire [0:1] mux_tree_tapbuf_size2_188_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_189_sram;
wire [0:1] mux_tree_tapbuf_size2_189_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_190_sram;
wire [0:1] mux_tree_tapbuf_size2_190_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_191_sram;
wire [0:1] mux_tree_tapbuf_size2_191_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_192_sram;
wire [0:1] mux_tree_tapbuf_size2_192_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_193_sram;
wire [0:1] mux_tree_tapbuf_size2_193_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_194_sram;
wire [0:1] mux_tree_tapbuf_size2_194_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_195_sram;
wire [0:1] mux_tree_tapbuf_size2_195_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_196_sram;
wire [0:1] mux_tree_tapbuf_size2_196_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_197_sram;
wire [0:1] mux_tree_tapbuf_size2_197_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_198_sram;
wire [0:1] mux_tree_tapbuf_size2_198_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_199_sram;
wire [0:1] mux_tree_tapbuf_size2_199_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_200_sram;
wire [0:1] mux_tree_tapbuf_size2_200_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_201_sram;
wire [0:1] mux_tree_tapbuf_size2_201_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_202_sram;
wire [0:1] mux_tree_tapbuf_size2_202_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_203_sram;
wire [0:1] mux_tree_tapbuf_size2_203_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_204_sram;
wire [0:1] mux_tree_tapbuf_size2_204_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_205_sram;
wire [0:1] mux_tree_tapbuf_size2_205_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_206_sram;
wire [0:1] mux_tree_tapbuf_size2_206_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_207_sram;
wire [0:1] mux_tree_tapbuf_size2_207_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_208_sram;
wire [0:1] mux_tree_tapbuf_size2_208_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_209_sram;
wire [0:1] mux_tree_tapbuf_size2_209_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_210_sram;
wire [0:1] mux_tree_tapbuf_size2_210_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_211_sram;
wire [0:1] mux_tree_tapbuf_size2_211_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_212_sram;
wire [0:1] mux_tree_tapbuf_size2_212_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_213_sram;
wire [0:1] mux_tree_tapbuf_size2_213_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_214_sram;
wire [0:1] mux_tree_tapbuf_size2_214_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_215_out;
wire [0:1] mux_tree_tapbuf_size2_215_sram;
wire [0:1] mux_tree_tapbuf_size2_215_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_216_out;
wire [0:1] mux_tree_tapbuf_size2_216_sram;
wire [0:1] mux_tree_tapbuf_size2_216_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_217_out;
wire [0:1] mux_tree_tapbuf_size2_217_sram;
wire [0:1] mux_tree_tapbuf_size2_217_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_218_out;
wire [0:1] mux_tree_tapbuf_size2_218_sram;
wire [0:1] mux_tree_tapbuf_size2_218_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_219_out;
wire [0:1] mux_tree_tapbuf_size2_219_sram;
wire [0:1] mux_tree_tapbuf_size2_219_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_220_out;
wire [0:1] mux_tree_tapbuf_size2_220_sram;
wire [0:1] mux_tree_tapbuf_size2_220_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_221_out;
wire [0:1] mux_tree_tapbuf_size2_221_sram;
wire [0:1] mux_tree_tapbuf_size2_221_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_222_out;
wire [0:1] mux_tree_tapbuf_size2_222_sram;
wire [0:1] mux_tree_tapbuf_size2_222_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_223_out;
wire [0:1] mux_tree_tapbuf_size2_223_sram;
wire [0:1] mux_tree_tapbuf_size2_223_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_224_out;
wire [0:1] mux_tree_tapbuf_size2_224_sram;
wire [0:1] mux_tree_tapbuf_size2_224_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_225_out;
wire [0:1] mux_tree_tapbuf_size2_225_sram;
wire [0:1] mux_tree_tapbuf_size2_225_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_226_out;
wire [0:1] mux_tree_tapbuf_size2_226_sram;
wire [0:1] mux_tree_tapbuf_size2_226_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_227_out;
wire [0:1] mux_tree_tapbuf_size2_227_sram;
wire [0:1] mux_tree_tapbuf_size2_227_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_228_out;
wire [0:1] mux_tree_tapbuf_size2_228_sram;
wire [0:1] mux_tree_tapbuf_size2_228_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_229_out;
wire [0:1] mux_tree_tapbuf_size2_229_sram;
wire [0:1] mux_tree_tapbuf_size2_229_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_230_out;
wire [0:1] mux_tree_tapbuf_size2_230_sram;
wire [0:1] mux_tree_tapbuf_size2_230_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_231_out;
wire [0:1] mux_tree_tapbuf_size2_231_sram;
wire [0:1] mux_tree_tapbuf_size2_231_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_232_out;
wire [0:1] mux_tree_tapbuf_size2_232_sram;
wire [0:1] mux_tree_tapbuf_size2_232_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_233_out;
wire [0:1] mux_tree_tapbuf_size2_233_sram;
wire [0:1] mux_tree_tapbuf_size2_233_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_234_out;
wire [0:1] mux_tree_tapbuf_size2_234_sram;
wire [0:1] mux_tree_tapbuf_size2_234_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_235_out;
wire [0:1] mux_tree_tapbuf_size2_235_sram;
wire [0:1] mux_tree_tapbuf_size2_235_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_236_out;
wire [0:1] mux_tree_tapbuf_size2_236_sram;
wire [0:1] mux_tree_tapbuf_size2_236_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_237_out;
wire [0:1] mux_tree_tapbuf_size2_237_sram;
wire [0:1] mux_tree_tapbuf_size2_237_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_238_out;
wire [0:1] mux_tree_tapbuf_size2_238_sram;
wire [0:1] mux_tree_tapbuf_size2_238_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_239_out;
wire [0:1] mux_tree_tapbuf_size2_239_sram;
wire [0:1] mux_tree_tapbuf_size2_239_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_240_out;
wire [0:1] mux_tree_tapbuf_size2_240_sram;
wire [0:1] mux_tree_tapbuf_size2_240_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_241_out;
wire [0:1] mux_tree_tapbuf_size2_241_sram;
wire [0:1] mux_tree_tapbuf_size2_241_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_242_out;
wire [0:1] mux_tree_tapbuf_size2_242_sram;
wire [0:1] mux_tree_tapbuf_size2_242_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_243_out;
wire [0:1] mux_tree_tapbuf_size2_243_sram;
wire [0:1] mux_tree_tapbuf_size2_243_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_244_out;
wire [0:1] mux_tree_tapbuf_size2_244_sram;
wire [0:1] mux_tree_tapbuf_size2_244_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_245_out;
wire [0:1] mux_tree_tapbuf_size2_245_sram;
wire [0:1] mux_tree_tapbuf_size2_245_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_246_out;
wire [0:1] mux_tree_tapbuf_size2_246_sram;
wire [0:1] mux_tree_tapbuf_size2_246_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_247_out;
wire [0:1] mux_tree_tapbuf_size2_247_sram;
wire [0:1] mux_tree_tapbuf_size2_247_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_248_out;
wire [0:1] mux_tree_tapbuf_size2_248_sram;
wire [0:1] mux_tree_tapbuf_size2_248_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_249_out;
wire [0:1] mux_tree_tapbuf_size2_249_sram;
wire [0:1] mux_tree_tapbuf_size2_249_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_250_out;
wire [0:1] mux_tree_tapbuf_size2_250_sram;
wire [0:1] mux_tree_tapbuf_size2_250_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_251_out;
wire [0:1] mux_tree_tapbuf_size2_251_sram;
wire [0:1] mux_tree_tapbuf_size2_251_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_252_out;
wire [0:1] mux_tree_tapbuf_size2_252_sram;
wire [0:1] mux_tree_tapbuf_size2_252_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_253_out;
wire [0:1] mux_tree_tapbuf_size2_253_sram;
wire [0:1] mux_tree_tapbuf_size2_253_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_254_out;
wire [0:1] mux_tree_tapbuf_size2_254_sram;
wire [0:1] mux_tree_tapbuf_size2_254_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_255_out;
wire [0:1] mux_tree_tapbuf_size2_255_sram;
wire [0:1] mux_tree_tapbuf_size2_255_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_256_out;
wire [0:1] mux_tree_tapbuf_size2_256_sram;
wire [0:1] mux_tree_tapbuf_size2_256_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_257_out;
wire [0:1] mux_tree_tapbuf_size2_257_sram;
wire [0:1] mux_tree_tapbuf_size2_257_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_258_out;
wire [0:1] mux_tree_tapbuf_size2_258_sram;
wire [0:1] mux_tree_tapbuf_size2_258_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_259_out;
wire [0:1] mux_tree_tapbuf_size2_259_sram;
wire [0:1] mux_tree_tapbuf_size2_259_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_260_out;
wire [0:1] mux_tree_tapbuf_size2_260_sram;
wire [0:1] mux_tree_tapbuf_size2_260_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_261_out;
wire [0:1] mux_tree_tapbuf_size2_261_sram;
wire [0:1] mux_tree_tapbuf_size2_261_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_262_out;
wire [0:1] mux_tree_tapbuf_size2_262_sram;
wire [0:1] mux_tree_tapbuf_size2_262_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_263_out;
wire [0:1] mux_tree_tapbuf_size2_263_sram;
wire [0:1] mux_tree_tapbuf_size2_263_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_264_out;
wire [0:1] mux_tree_tapbuf_size2_264_sram;
wire [0:1] mux_tree_tapbuf_size2_264_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_265_out;
wire [0:1] mux_tree_tapbuf_size2_265_sram;
wire [0:1] mux_tree_tapbuf_size2_265_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_266_out;
wire [0:1] mux_tree_tapbuf_size2_266_sram;
wire [0:1] mux_tree_tapbuf_size2_266_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_267_out;
wire [0:1] mux_tree_tapbuf_size2_267_sram;
wire [0:1] mux_tree_tapbuf_size2_267_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_268_out;
wire [0:1] mux_tree_tapbuf_size2_268_sram;
wire [0:1] mux_tree_tapbuf_size2_268_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_269_out;
wire [0:1] mux_tree_tapbuf_size2_269_sram;
wire [0:1] mux_tree_tapbuf_size2_269_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_270_out;
wire [0:1] mux_tree_tapbuf_size2_270_sram;
wire [0:1] mux_tree_tapbuf_size2_270_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_271_out;
wire [0:1] mux_tree_tapbuf_size2_271_sram;
wire [0:1] mux_tree_tapbuf_size2_271_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_272_out;
wire [0:1] mux_tree_tapbuf_size2_272_sram;
wire [0:1] mux_tree_tapbuf_size2_272_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_273_out;
wire [0:1] mux_tree_tapbuf_size2_273_sram;
wire [0:1] mux_tree_tapbuf_size2_273_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_274_out;
wire [0:1] mux_tree_tapbuf_size2_274_sram;
wire [0:1] mux_tree_tapbuf_size2_274_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_275_out;
wire [0:1] mux_tree_tapbuf_size2_275_sram;
wire [0:1] mux_tree_tapbuf_size2_275_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_276_out;
wire [0:1] mux_tree_tapbuf_size2_276_sram;
wire [0:1] mux_tree_tapbuf_size2_276_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_277_out;
wire [0:1] mux_tree_tapbuf_size2_277_sram;
wire [0:1] mux_tree_tapbuf_size2_277_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_278_out;
wire [0:1] mux_tree_tapbuf_size2_278_sram;
wire [0:1] mux_tree_tapbuf_size2_278_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_279_out;
wire [0:1] mux_tree_tapbuf_size2_279_sram;
wire [0:1] mux_tree_tapbuf_size2_279_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_280_out;
wire [0:1] mux_tree_tapbuf_size2_280_sram;
wire [0:1] mux_tree_tapbuf_size2_280_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_281_out;
wire [0:1] mux_tree_tapbuf_size2_281_sram;
wire [0:1] mux_tree_tapbuf_size2_281_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_282_out;
wire [0:1] mux_tree_tapbuf_size2_282_sram;
wire [0:1] mux_tree_tapbuf_size2_282_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_283_out;
wire [0:1] mux_tree_tapbuf_size2_283_sram;
wire [0:1] mux_tree_tapbuf_size2_283_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_284_out;
wire [0:1] mux_tree_tapbuf_size2_284_sram;
wire [0:1] mux_tree_tapbuf_size2_284_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_285_out;
wire [0:1] mux_tree_tapbuf_size2_285_sram;
wire [0:1] mux_tree_tapbuf_size2_285_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_286_out;
wire [0:1] mux_tree_tapbuf_size2_286_sram;
wire [0:1] mux_tree_tapbuf_size2_286_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_287_out;
wire [0:1] mux_tree_tapbuf_size2_287_sram;
wire [0:1] mux_tree_tapbuf_size2_287_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_288_out;
wire [0:1] mux_tree_tapbuf_size2_288_sram;
wire [0:1] mux_tree_tapbuf_size2_288_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_289_out;
wire [0:1] mux_tree_tapbuf_size2_289_sram;
wire [0:1] mux_tree_tapbuf_size2_289_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_290_out;
wire [0:1] mux_tree_tapbuf_size2_290_sram;
wire [0:1] mux_tree_tapbuf_size2_290_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_291_out;
wire [0:1] mux_tree_tapbuf_size2_291_sram;
wire [0:1] mux_tree_tapbuf_size2_291_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_292_out;
wire [0:1] mux_tree_tapbuf_size2_292_sram;
wire [0:1] mux_tree_tapbuf_size2_292_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_293_out;
wire [0:1] mux_tree_tapbuf_size2_293_sram;
wire [0:1] mux_tree_tapbuf_size2_293_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_294_out;
wire [0:1] mux_tree_tapbuf_size2_294_sram;
wire [0:1] mux_tree_tapbuf_size2_294_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_295_out;
wire [0:1] mux_tree_tapbuf_size2_295_sram;
wire [0:1] mux_tree_tapbuf_size2_295_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_296_out;
wire [0:1] mux_tree_tapbuf_size2_296_sram;
wire [0:1] mux_tree_tapbuf_size2_296_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_297_out;
wire [0:1] mux_tree_tapbuf_size2_297_sram;
wire [0:1] mux_tree_tapbuf_size2_297_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_298_out;
wire [0:1] mux_tree_tapbuf_size2_298_sram;
wire [0:1] mux_tree_tapbuf_size2_298_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_299_out;
wire [0:1] mux_tree_tapbuf_size2_299_sram;
wire [0:1] mux_tree_tapbuf_size2_299_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_300_out;
wire [0:1] mux_tree_tapbuf_size2_300_sram;
wire [0:1] mux_tree_tapbuf_size2_300_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_301_out;
wire [0:1] mux_tree_tapbuf_size2_301_sram;
wire [0:1] mux_tree_tapbuf_size2_301_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_302_out;
wire [0:1] mux_tree_tapbuf_size2_302_sram;
wire [0:1] mux_tree_tapbuf_size2_302_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_303_out;
wire [0:1] mux_tree_tapbuf_size2_303_sram;
wire [0:1] mux_tree_tapbuf_size2_303_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_304_out;
wire [0:1] mux_tree_tapbuf_size2_304_sram;
wire [0:1] mux_tree_tapbuf_size2_304_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_305_out;
wire [0:1] mux_tree_tapbuf_size2_305_sram;
wire [0:1] mux_tree_tapbuf_size2_305_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_306_out;
wire [0:1] mux_tree_tapbuf_size2_306_sram;
wire [0:1] mux_tree_tapbuf_size2_306_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_307_out;
wire [0:1] mux_tree_tapbuf_size2_307_sram;
wire [0:1] mux_tree_tapbuf_size2_307_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_308_out;
wire [0:1] mux_tree_tapbuf_size2_308_sram;
wire [0:1] mux_tree_tapbuf_size2_308_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_309_out;
wire [0:1] mux_tree_tapbuf_size2_309_sram;
wire [0:1] mux_tree_tapbuf_size2_309_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_310_out;
wire [0:1] mux_tree_tapbuf_size2_310_sram;
wire [0:1] mux_tree_tapbuf_size2_310_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_311_out;
wire [0:1] mux_tree_tapbuf_size2_311_sram;
wire [0:1] mux_tree_tapbuf_size2_311_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_312_out;
wire [0:1] mux_tree_tapbuf_size2_312_sram;
wire [0:1] mux_tree_tapbuf_size2_312_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_313_out;
wire [0:1] mux_tree_tapbuf_size2_313_sram;
wire [0:1] mux_tree_tapbuf_size2_313_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_314_out;
wire [0:1] mux_tree_tapbuf_size2_314_sram;
wire [0:1] mux_tree_tapbuf_size2_314_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_315_out;
wire [0:1] mux_tree_tapbuf_size2_315_sram;
wire [0:1] mux_tree_tapbuf_size2_315_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_316_out;
wire [0:1] mux_tree_tapbuf_size2_316_sram;
wire [0:1] mux_tree_tapbuf_size2_316_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_317_out;
wire [0:1] mux_tree_tapbuf_size2_317_sram;
wire [0:1] mux_tree_tapbuf_size2_317_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_318_out;
wire [0:1] mux_tree_tapbuf_size2_318_sram;
wire [0:1] mux_tree_tapbuf_size2_318_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_319_out;
wire [0:1] mux_tree_tapbuf_size2_319_sram;
wire [0:1] mux_tree_tapbuf_size2_319_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_320_out;
wire [0:1] mux_tree_tapbuf_size2_320_sram;
wire [0:1] mux_tree_tapbuf_size2_320_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_321_out;
wire [0:1] mux_tree_tapbuf_size2_321_sram;
wire [0:1] mux_tree_tapbuf_size2_321_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_322_out;
wire [0:1] mux_tree_tapbuf_size2_322_sram;
wire [0:1] mux_tree_tapbuf_size2_322_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_323_out;
wire [0:1] mux_tree_tapbuf_size2_323_sram;
wire [0:1] mux_tree_tapbuf_size2_323_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_324_out;
wire [0:1] mux_tree_tapbuf_size2_324_sram;
wire [0:1] mux_tree_tapbuf_size2_324_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_325_out;
wire [0:1] mux_tree_tapbuf_size2_325_sram;
wire [0:1] mux_tree_tapbuf_size2_325_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_326_out;
wire [0:1] mux_tree_tapbuf_size2_326_sram;
wire [0:1] mux_tree_tapbuf_size2_326_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_327_out;
wire [0:1] mux_tree_tapbuf_size2_327_sram;
wire [0:1] mux_tree_tapbuf_size2_327_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_328_out;
wire [0:1] mux_tree_tapbuf_size2_328_sram;
wire [0:1] mux_tree_tapbuf_size2_328_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_329_out;
wire [0:1] mux_tree_tapbuf_size2_329_sram;
wire [0:1] mux_tree_tapbuf_size2_329_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_330_out;
wire [0:1] mux_tree_tapbuf_size2_330_sram;
wire [0:1] mux_tree_tapbuf_size2_330_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_331_out;
wire [0:1] mux_tree_tapbuf_size2_331_sram;
wire [0:1] mux_tree_tapbuf_size2_331_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_332_out;
wire [0:1] mux_tree_tapbuf_size2_332_sram;
wire [0:1] mux_tree_tapbuf_size2_332_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_333_out;
wire [0:1] mux_tree_tapbuf_size2_333_sram;
wire [0:1] mux_tree_tapbuf_size2_333_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_334_out;
wire [0:1] mux_tree_tapbuf_size2_334_sram;
wire [0:1] mux_tree_tapbuf_size2_334_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_335_out;
wire [0:1] mux_tree_tapbuf_size2_335_sram;
wire [0:1] mux_tree_tapbuf_size2_335_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_336_out;
wire [0:1] mux_tree_tapbuf_size2_336_sram;
wire [0:1] mux_tree_tapbuf_size2_336_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_337_out;
wire [0:1] mux_tree_tapbuf_size2_337_sram;
wire [0:1] mux_tree_tapbuf_size2_337_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_338_out;
wire [0:1] mux_tree_tapbuf_size2_338_sram;
wire [0:1] mux_tree_tapbuf_size2_338_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_339_out;
wire [0:1] mux_tree_tapbuf_size2_339_sram;
wire [0:1] mux_tree_tapbuf_size2_339_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_340_out;
wire [0:1] mux_tree_tapbuf_size2_340_sram;
wire [0:1] mux_tree_tapbuf_size2_340_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_341_out;
wire [0:1] mux_tree_tapbuf_size2_341_sram;
wire [0:1] mux_tree_tapbuf_size2_341_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_342_out;
wire [0:1] mux_tree_tapbuf_size2_342_sram;
wire [0:1] mux_tree_tapbuf_size2_342_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_343_out;
wire [0:1] mux_tree_tapbuf_size2_343_sram;
wire [0:1] mux_tree_tapbuf_size2_343_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_344_out;
wire [0:1] mux_tree_tapbuf_size2_344_sram;
wire [0:1] mux_tree_tapbuf_size2_344_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_345_out;
wire [0:1] mux_tree_tapbuf_size2_345_sram;
wire [0:1] mux_tree_tapbuf_size2_345_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_346_out;
wire [0:1] mux_tree_tapbuf_size2_346_sram;
wire [0:1] mux_tree_tapbuf_size2_346_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_347_out;
wire [0:1] mux_tree_tapbuf_size2_347_sram;
wire [0:1] mux_tree_tapbuf_size2_347_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_348_out;
wire [0:1] mux_tree_tapbuf_size2_348_sram;
wire [0:1] mux_tree_tapbuf_size2_348_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_349_out;
wire [0:1] mux_tree_tapbuf_size2_349_sram;
wire [0:1] mux_tree_tapbuf_size2_349_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_350_out;
wire [0:1] mux_tree_tapbuf_size2_350_sram;
wire [0:1] mux_tree_tapbuf_size2_350_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_351_out;
wire [0:1] mux_tree_tapbuf_size2_351_sram;
wire [0:1] mux_tree_tapbuf_size2_351_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_352_out;
wire [0:1] mux_tree_tapbuf_size2_352_sram;
wire [0:1] mux_tree_tapbuf_size2_352_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_353_out;
wire [0:1] mux_tree_tapbuf_size2_353_sram;
wire [0:1] mux_tree_tapbuf_size2_353_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_354_out;
wire [0:1] mux_tree_tapbuf_size2_354_sram;
wire [0:1] mux_tree_tapbuf_size2_354_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_355_out;
wire [0:1] mux_tree_tapbuf_size2_355_sram;
wire [0:1] mux_tree_tapbuf_size2_355_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_356_out;
wire [0:1] mux_tree_tapbuf_size2_356_sram;
wire [0:1] mux_tree_tapbuf_size2_356_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_357_out;
wire [0:1] mux_tree_tapbuf_size2_357_sram;
wire [0:1] mux_tree_tapbuf_size2_357_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_358_out;
wire [0:1] mux_tree_tapbuf_size2_358_sram;
wire [0:1] mux_tree_tapbuf_size2_358_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_359_out;
wire [0:1] mux_tree_tapbuf_size2_359_sram;
wire [0:1] mux_tree_tapbuf_size2_359_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_360_out;
wire [0:1] mux_tree_tapbuf_size2_360_sram;
wire [0:1] mux_tree_tapbuf_size2_360_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_361_out;
wire [0:1] mux_tree_tapbuf_size2_361_sram;
wire [0:1] mux_tree_tapbuf_size2_361_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_362_out;
wire [0:1] mux_tree_tapbuf_size2_362_sram;
wire [0:1] mux_tree_tapbuf_size2_362_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_363_out;
wire [0:1] mux_tree_tapbuf_size2_363_sram;
wire [0:1] mux_tree_tapbuf_size2_363_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_364_out;
wire [0:1] mux_tree_tapbuf_size2_364_sram;
wire [0:1] mux_tree_tapbuf_size2_364_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_365_out;
wire [0:1] mux_tree_tapbuf_size2_365_sram;
wire [0:1] mux_tree_tapbuf_size2_365_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_366_out;
wire [0:1] mux_tree_tapbuf_size2_366_sram;
wire [0:1] mux_tree_tapbuf_size2_366_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_367_out;
wire [0:1] mux_tree_tapbuf_size2_367_sram;
wire [0:1] mux_tree_tapbuf_size2_367_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_368_out;
wire [0:1] mux_tree_tapbuf_size2_368_sram;
wire [0:1] mux_tree_tapbuf_size2_368_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_369_out;
wire [0:1] mux_tree_tapbuf_size2_369_sram;
wire [0:1] mux_tree_tapbuf_size2_369_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_370_out;
wire [0:1] mux_tree_tapbuf_size2_370_sram;
wire [0:1] mux_tree_tapbuf_size2_370_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_371_out;
wire [0:1] mux_tree_tapbuf_size2_371_sram;
wire [0:1] mux_tree_tapbuf_size2_371_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_372_out;
wire [0:1] mux_tree_tapbuf_size2_372_sram;
wire [0:1] mux_tree_tapbuf_size2_372_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_373_out;
wire [0:1] mux_tree_tapbuf_size2_373_sram;
wire [0:1] mux_tree_tapbuf_size2_373_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_374_out;
wire [0:1] mux_tree_tapbuf_size2_374_sram;
wire [0:1] mux_tree_tapbuf_size2_374_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_375_out;
wire [0:1] mux_tree_tapbuf_size2_375_sram;
wire [0:1] mux_tree_tapbuf_size2_375_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_376_out;
wire [0:1] mux_tree_tapbuf_size2_376_sram;
wire [0:1] mux_tree_tapbuf_size2_376_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_377_out;
wire [0:1] mux_tree_tapbuf_size2_377_sram;
wire [0:1] mux_tree_tapbuf_size2_377_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_378_out;
wire [0:1] mux_tree_tapbuf_size2_378_sram;
wire [0:1] mux_tree_tapbuf_size2_378_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_379_out;
wire [0:1] mux_tree_tapbuf_size2_379_sram;
wire [0:1] mux_tree_tapbuf_size2_379_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_380_out;
wire [0:1] mux_tree_tapbuf_size2_380_sram;
wire [0:1] mux_tree_tapbuf_size2_380_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_381_out;
wire [0:1] mux_tree_tapbuf_size2_381_sram;
wire [0:1] mux_tree_tapbuf_size2_381_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_382_out;
wire [0:1] mux_tree_tapbuf_size2_382_sram;
wire [0:1] mux_tree_tapbuf_size2_382_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_383_out;
wire [0:1] mux_tree_tapbuf_size2_383_sram;
wire [0:1] mux_tree_tapbuf_size2_383_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_384_out;
wire [0:1] mux_tree_tapbuf_size2_384_sram;
wire [0:1] mux_tree_tapbuf_size2_384_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_385_out;
wire [0:1] mux_tree_tapbuf_size2_385_sram;
wire [0:1] mux_tree_tapbuf_size2_385_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_386_out;
wire [0:1] mux_tree_tapbuf_size2_386_sram;
wire [0:1] mux_tree_tapbuf_size2_386_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_387_out;
wire [0:1] mux_tree_tapbuf_size2_387_sram;
wire [0:1] mux_tree_tapbuf_size2_387_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_388_out;
wire [0:1] mux_tree_tapbuf_size2_388_sram;
wire [0:1] mux_tree_tapbuf_size2_388_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_389_out;
wire [0:1] mux_tree_tapbuf_size2_389_sram;
wire [0:1] mux_tree_tapbuf_size2_389_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_390_out;
wire [0:1] mux_tree_tapbuf_size2_390_sram;
wire [0:1] mux_tree_tapbuf_size2_390_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_391_out;
wire [0:1] mux_tree_tapbuf_size2_391_sram;
wire [0:1] mux_tree_tapbuf_size2_391_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_392_out;
wire [0:1] mux_tree_tapbuf_size2_392_sram;
wire [0:1] mux_tree_tapbuf_size2_392_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_393_out;
wire [0:1] mux_tree_tapbuf_size2_393_sram;
wire [0:1] mux_tree_tapbuf_size2_393_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_394_out;
wire [0:1] mux_tree_tapbuf_size2_394_sram;
wire [0:1] mux_tree_tapbuf_size2_394_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_395_out;
wire [0:1] mux_tree_tapbuf_size2_395_sram;
wire [0:1] mux_tree_tapbuf_size2_395_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_396_out;
wire [0:1] mux_tree_tapbuf_size2_396_sram;
wire [0:1] mux_tree_tapbuf_size2_396_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_397_out;
wire [0:1] mux_tree_tapbuf_size2_397_sram;
wire [0:1] mux_tree_tapbuf_size2_397_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_398_out;
wire [0:1] mux_tree_tapbuf_size2_398_sram;
wire [0:1] mux_tree_tapbuf_size2_398_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_399_out;
wire [0:1] mux_tree_tapbuf_size2_399_sram;
wire [0:1] mux_tree_tapbuf_size2_399_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_400_out;
wire [0:1] mux_tree_tapbuf_size2_400_sram;
wire [0:1] mux_tree_tapbuf_size2_400_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_401_out;
wire [0:1] mux_tree_tapbuf_size2_401_sram;
wire [0:1] mux_tree_tapbuf_size2_401_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_402_out;
wire [0:1] mux_tree_tapbuf_size2_402_sram;
wire [0:1] mux_tree_tapbuf_size2_402_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_403_out;
wire [0:1] mux_tree_tapbuf_size2_403_sram;
wire [0:1] mux_tree_tapbuf_size2_403_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_404_out;
wire [0:1] mux_tree_tapbuf_size2_404_sram;
wire [0:1] mux_tree_tapbuf_size2_404_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_405_out;
wire [0:1] mux_tree_tapbuf_size2_405_sram;
wire [0:1] mux_tree_tapbuf_size2_405_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_406_out;
wire [0:1] mux_tree_tapbuf_size2_406_sram;
wire [0:1] mux_tree_tapbuf_size2_406_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_407_out;
wire [0:1] mux_tree_tapbuf_size2_407_sram;
wire [0:1] mux_tree_tapbuf_size2_407_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_408_out;
wire [0:1] mux_tree_tapbuf_size2_408_sram;
wire [0:1] mux_tree_tapbuf_size2_408_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_409_out;
wire [0:1] mux_tree_tapbuf_size2_409_sram;
wire [0:1] mux_tree_tapbuf_size2_409_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_40_sram;
wire [0:1] mux_tree_tapbuf_size2_40_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_410_out;
wire [0:1] mux_tree_tapbuf_size2_410_sram;
wire [0:1] mux_tree_tapbuf_size2_410_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_411_out;
wire [0:1] mux_tree_tapbuf_size2_411_sram;
wire [0:1] mux_tree_tapbuf_size2_411_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_412_out;
wire [0:1] mux_tree_tapbuf_size2_412_sram;
wire [0:1] mux_tree_tapbuf_size2_412_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_413_out;
wire [0:1] mux_tree_tapbuf_size2_413_sram;
wire [0:1] mux_tree_tapbuf_size2_413_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_414_out;
wire [0:1] mux_tree_tapbuf_size2_414_sram;
wire [0:1] mux_tree_tapbuf_size2_414_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_415_out;
wire [0:1] mux_tree_tapbuf_size2_415_sram;
wire [0:1] mux_tree_tapbuf_size2_415_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_416_out;
wire [0:1] mux_tree_tapbuf_size2_416_sram;
wire [0:1] mux_tree_tapbuf_size2_416_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_417_out;
wire [0:1] mux_tree_tapbuf_size2_417_sram;
wire [0:1] mux_tree_tapbuf_size2_417_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_418_out;
wire [0:1] mux_tree_tapbuf_size2_418_sram;
wire [0:1] mux_tree_tapbuf_size2_418_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_419_out;
wire [0:1] mux_tree_tapbuf_size2_419_sram;
wire [0:1] mux_tree_tapbuf_size2_419_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_41_sram;
wire [0:1] mux_tree_tapbuf_size2_41_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_420_out;
wire [0:1] mux_tree_tapbuf_size2_420_sram;
wire [0:1] mux_tree_tapbuf_size2_420_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_421_out;
wire [0:1] mux_tree_tapbuf_size2_421_sram;
wire [0:1] mux_tree_tapbuf_size2_421_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_422_out;
wire [0:1] mux_tree_tapbuf_size2_422_sram;
wire [0:1] mux_tree_tapbuf_size2_422_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_423_out;
wire [0:1] mux_tree_tapbuf_size2_423_sram;
wire [0:1] mux_tree_tapbuf_size2_423_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_424_out;
wire [0:1] mux_tree_tapbuf_size2_424_sram;
wire [0:1] mux_tree_tapbuf_size2_424_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_42_sram;
wire [0:1] mux_tree_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_43_sram;
wire [0:1] mux_tree_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_44_sram;
wire [0:1] mux_tree_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_45_sram;
wire [0:1] mux_tree_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_46_sram;
wire [0:1] mux_tree_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_47_sram;
wire [0:1] mux_tree_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_48_sram;
wire [0:1] mux_tree_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_49_sram;
wire [0:1] mux_tree_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_50_sram;
wire [0:1] mux_tree_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_51_sram;
wire [0:1] mux_tree_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_52_sram;
wire [0:1] mux_tree_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_53_sram;
wire [0:1] mux_tree_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_54_sram;
wire [0:1] mux_tree_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_55_sram;
wire [0:1] mux_tree_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_56_sram;
wire [0:1] mux_tree_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_57_sram;
wire [0:1] mux_tree_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_58_sram;
wire [0:1] mux_tree_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_59_sram;
wire [0:1] mux_tree_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_60_sram;
wire [0:1] mux_tree_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_61_sram;
wire [0:1] mux_tree_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_62_sram;
wire [0:1] mux_tree_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_63_sram;
wire [0:1] mux_tree_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_64_sram;
wire [0:1] mux_tree_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_65_sram;
wire [0:1] mux_tree_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_66_sram;
wire [0:1] mux_tree_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_67_sram;
wire [0:1] mux_tree_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_68_sram;
wire [0:1] mux_tree_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_69_sram;
wire [0:1] mux_tree_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_70_sram;
wire [0:1] mux_tree_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_71_sram;
wire [0:1] mux_tree_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_72_sram;
wire [0:1] mux_tree_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_73_sram;
wire [0:1] mux_tree_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_74_sram;
wire [0:1] mux_tree_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_75_sram;
wire [0:1] mux_tree_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_76_sram;
wire [0:1] mux_tree_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_77_sram;
wire [0:1] mux_tree_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_78_sram;
wire [0:1] mux_tree_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_79_sram;
wire [0:1] mux_tree_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_80_sram;
wire [0:1] mux_tree_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_81_sram;
wire [0:1] mux_tree_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_82_sram;
wire [0:1] mux_tree_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_83_sram;
wire [0:1] mux_tree_tapbuf_size2_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_84_sram;
wire [0:1] mux_tree_tapbuf_size2_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_85_sram;
wire [0:1] mux_tree_tapbuf_size2_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_86_sram;
wire [0:1] mux_tree_tapbuf_size2_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_87_sram;
wire [0:1] mux_tree_tapbuf_size2_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_88_sram;
wire [0:1] mux_tree_tapbuf_size2_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_89_sram;
wire [0:1] mux_tree_tapbuf_size2_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_90_sram;
wire [0:1] mux_tree_tapbuf_size2_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_91_sram;
wire [0:1] mux_tree_tapbuf_size2_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_92_sram;
wire [0:1] mux_tree_tapbuf_size2_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_93_sram;
wire [0:1] mux_tree_tapbuf_size2_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_94_sram;
wire [0:1] mux_tree_tapbuf_size2_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_95_sram;
wire [0:1] mux_tree_tapbuf_size2_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_96_sram;
wire [0:1] mux_tree_tapbuf_size2_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_97_sram;
wire [0:1] mux_tree_tapbuf_size2_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_98_sram;
wire [0:1] mux_tree_tapbuf_size2_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_99_sram;
wire [0:1] mux_tree_tapbuf_size2_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_225_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_226_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_227_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_228_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_229_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_230_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_231_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_232_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_233_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_234_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_235_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_236_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_237_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_238_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_239_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_240_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_241_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_242_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_243_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_244_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_245_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_246_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_247_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_248_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_249_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_250_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_251_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_252_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_253_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_254_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_255_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_256_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_257_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_258_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_259_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_260_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_261_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_262_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_263_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_264_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_265_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_266_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_267_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_268_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_269_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_270_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_271_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_272_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_273_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_274_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_275_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_276_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_277_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_278_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_279_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_280_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_281_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_282_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_283_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_284_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_285_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_286_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_287_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_288_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_289_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_290_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_291_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_292_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_293_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_294_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_295_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_296_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_297_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_298_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_299_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_300_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_301_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_302_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_303_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_304_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_305_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_306_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_307_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_308_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_309_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_310_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_311_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_312_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_313_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_314_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_315_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_316_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_317_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_318_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_319_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_320_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_321_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_322_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_323_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_324_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_325_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_326_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_327_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_328_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_329_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_330_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_331_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_332_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_333_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_334_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_335_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_336_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_337_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_338_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_339_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_340_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_341_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_342_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_343_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_344_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_345_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_346_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_347_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_348_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_349_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_350_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_351_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_352_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_353_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_354_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_355_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_356_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_357_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_358_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_359_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_360_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_361_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_362_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_363_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_364_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_365_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_366_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_367_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_368_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_369_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_370_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_371_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_372_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_373_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_374_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_375_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_376_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_377_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_378_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_379_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_380_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_381_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_382_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_383_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_384_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_385_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_386_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_387_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_388_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_389_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_390_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_391_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_392_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_393_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_394_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_395_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_396_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_397_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_398_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_399_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_400_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_401_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_402_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_403_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_404_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_405_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_406_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_407_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_408_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_409_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_410_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_411_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_412_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_413_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_414_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_415_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_416_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_417_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_418_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_419_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_420_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_421_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_422_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_423_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0 (
		.clk(clk),
		.router_wrap_RST_(mux_tree_tapbuf_size2_215_out),
		.router_wrap_MY_XPOS({mux_tree_tapbuf_size2_216_out, mux_tree_tapbuf_size2_217_out}),
		.router_wrap_MY_YPOS({mux_tree_tapbuf_size2_218_out, mux_tree_tapbuf_size2_219_out}),
		.router_wrap_IDATA_0({mux_tree_tapbuf_size2_220_out, mux_tree_tapbuf_size2_221_out, mux_tree_tapbuf_size2_222_out, mux_tree_tapbuf_size2_223_out, mux_tree_tapbuf_size2_224_out, mux_tree_tapbuf_size2_225_out, mux_tree_tapbuf_size2_226_out, mux_tree_tapbuf_size2_227_out, mux_tree_tapbuf_size2_228_out, mux_tree_tapbuf_size2_229_out, mux_tree_tapbuf_size2_230_out, mux_tree_tapbuf_size2_231_out, mux_tree_tapbuf_size2_232_out, mux_tree_tapbuf_size2_233_out, mux_tree_tapbuf_size2_234_out, mux_tree_tapbuf_size2_235_out, mux_tree_tapbuf_size2_236_out, mux_tree_tapbuf_size2_237_out, mux_tree_tapbuf_size2_238_out, mux_tree_tapbuf_size2_239_out, mux_tree_tapbuf_size2_240_out, mux_tree_tapbuf_size2_241_out, mux_tree_tapbuf_size2_242_out, mux_tree_tapbuf_size2_243_out, mux_tree_tapbuf_size2_244_out, mux_tree_tapbuf_size2_245_out, mux_tree_tapbuf_size2_246_out, mux_tree_tapbuf_size2_247_out, mux_tree_tapbuf_size2_248_out, mux_tree_tapbuf_size2_249_out, mux_tree_tapbuf_size2_250_out, mux_tree_tapbuf_size2_251_out, mux_tree_tapbuf_size2_252_out, mux_tree_tapbuf_size2_253_out, mux_tree_tapbuf_size2_254_out}),
		.router_wrap_IDATA_1({mux_tree_tapbuf_size2_255_out, mux_tree_tapbuf_size2_256_out, mux_tree_tapbuf_size2_257_out, mux_tree_tapbuf_size2_258_out, mux_tree_tapbuf_size2_259_out, mux_tree_tapbuf_size2_260_out, mux_tree_tapbuf_size2_261_out, mux_tree_tapbuf_size2_262_out, mux_tree_tapbuf_size2_263_out, mux_tree_tapbuf_size2_264_out, mux_tree_tapbuf_size2_265_out, mux_tree_tapbuf_size2_266_out, mux_tree_tapbuf_size2_267_out, mux_tree_tapbuf_size2_268_out, mux_tree_tapbuf_size2_269_out, mux_tree_tapbuf_size2_270_out, mux_tree_tapbuf_size2_271_out, mux_tree_tapbuf_size2_272_out, mux_tree_tapbuf_size2_273_out, mux_tree_tapbuf_size2_274_out, mux_tree_tapbuf_size2_275_out, mux_tree_tapbuf_size2_276_out, mux_tree_tapbuf_size2_277_out, mux_tree_tapbuf_size2_278_out, mux_tree_tapbuf_size2_279_out, mux_tree_tapbuf_size2_280_out, mux_tree_tapbuf_size2_281_out, mux_tree_tapbuf_size2_282_out, mux_tree_tapbuf_size2_283_out, mux_tree_tapbuf_size2_284_out, mux_tree_tapbuf_size2_285_out, mux_tree_tapbuf_size2_286_out, mux_tree_tapbuf_size2_287_out, mux_tree_tapbuf_size2_288_out, mux_tree_tapbuf_size2_289_out}),
		.router_wrap_IDATA_2({mux_tree_tapbuf_size2_290_out, mux_tree_tapbuf_size2_291_out, mux_tree_tapbuf_size2_292_out, mux_tree_tapbuf_size2_293_out, mux_tree_tapbuf_size2_294_out, mux_tree_tapbuf_size2_295_out, mux_tree_tapbuf_size2_296_out, mux_tree_tapbuf_size2_297_out, mux_tree_tapbuf_size2_298_out, mux_tree_tapbuf_size2_299_out, mux_tree_tapbuf_size2_300_out, mux_tree_tapbuf_size2_301_out, mux_tree_tapbuf_size2_302_out, mux_tree_tapbuf_size2_303_out, mux_tree_tapbuf_size2_304_out, mux_tree_tapbuf_size2_305_out, mux_tree_tapbuf_size2_306_out, mux_tree_tapbuf_size2_307_out, mux_tree_tapbuf_size2_308_out, mux_tree_tapbuf_size2_309_out, mux_tree_tapbuf_size2_310_out, mux_tree_tapbuf_size2_311_out, mux_tree_tapbuf_size2_312_out, mux_tree_tapbuf_size2_313_out, mux_tree_tapbuf_size2_314_out, mux_tree_tapbuf_size2_315_out, mux_tree_tapbuf_size2_316_out, mux_tree_tapbuf_size2_317_out, mux_tree_tapbuf_size2_318_out, mux_tree_tapbuf_size2_319_out, mux_tree_tapbuf_size2_320_out, mux_tree_tapbuf_size2_321_out, mux_tree_tapbuf_size2_322_out, mux_tree_tapbuf_size2_323_out, mux_tree_tapbuf_size2_324_out}),
		.router_wrap_IDATA_3({mux_tree_tapbuf_size2_325_out, mux_tree_tapbuf_size2_326_out, mux_tree_tapbuf_size2_327_out, mux_tree_tapbuf_size2_328_out, mux_tree_tapbuf_size2_329_out, mux_tree_tapbuf_size2_330_out, mux_tree_tapbuf_size2_331_out, mux_tree_tapbuf_size2_332_out, mux_tree_tapbuf_size2_333_out, mux_tree_tapbuf_size2_334_out, mux_tree_tapbuf_size2_335_out, mux_tree_tapbuf_size2_336_out, mux_tree_tapbuf_size2_337_out, mux_tree_tapbuf_size2_338_out, mux_tree_tapbuf_size2_339_out, mux_tree_tapbuf_size2_340_out, mux_tree_tapbuf_size2_341_out, mux_tree_tapbuf_size2_342_out, mux_tree_tapbuf_size2_343_out, mux_tree_tapbuf_size2_344_out, mux_tree_tapbuf_size2_345_out, mux_tree_tapbuf_size2_346_out, mux_tree_tapbuf_size2_347_out, mux_tree_tapbuf_size2_348_out, mux_tree_tapbuf_size2_349_out, mux_tree_tapbuf_size2_350_out, mux_tree_tapbuf_size2_351_out, mux_tree_tapbuf_size2_352_out, mux_tree_tapbuf_size2_353_out, mux_tree_tapbuf_size2_354_out, mux_tree_tapbuf_size2_355_out, mux_tree_tapbuf_size2_356_out, mux_tree_tapbuf_size2_357_out, mux_tree_tapbuf_size2_358_out, mux_tree_tapbuf_size2_359_out}),
		.router_wrap_IDATA_4({mux_tree_tapbuf_size2_360_out, mux_tree_tapbuf_size2_361_out, mux_tree_tapbuf_size2_362_out, mux_tree_tapbuf_size2_363_out, mux_tree_tapbuf_size2_364_out, mux_tree_tapbuf_size2_365_out, mux_tree_tapbuf_size2_366_out, mux_tree_tapbuf_size2_367_out, mux_tree_tapbuf_size2_368_out, mux_tree_tapbuf_size2_369_out, mux_tree_tapbuf_size2_370_out, mux_tree_tapbuf_size2_371_out, mux_tree_tapbuf_size2_372_out, mux_tree_tapbuf_size2_373_out, mux_tree_tapbuf_size2_374_out, mux_tree_tapbuf_size2_375_out, mux_tree_tapbuf_size2_376_out, mux_tree_tapbuf_size2_377_out, mux_tree_tapbuf_size2_378_out, mux_tree_tapbuf_size2_379_out, mux_tree_tapbuf_size2_380_out, mux_tree_tapbuf_size2_381_out, mux_tree_tapbuf_size2_382_out, mux_tree_tapbuf_size2_383_out, mux_tree_tapbuf_size2_384_out, mux_tree_tapbuf_size2_385_out, mux_tree_tapbuf_size2_386_out, mux_tree_tapbuf_size2_387_out, mux_tree_tapbuf_size2_388_out, mux_tree_tapbuf_size2_389_out, mux_tree_tapbuf_size2_390_out, mux_tree_tapbuf_size2_391_out, mux_tree_tapbuf_size2_392_out, mux_tree_tapbuf_size2_393_out, mux_tree_tapbuf_size2_394_out}),
		.router_wrap_IVALID_0(mux_tree_tapbuf_size2_395_out),
		.router_wrap_IVALID_1(mux_tree_tapbuf_size2_396_out),
		.router_wrap_IVALID_2(mux_tree_tapbuf_size2_397_out),
		.router_wrap_IVALID_3(mux_tree_tapbuf_size2_398_out),
		.router_wrap_IVALID_4(mux_tree_tapbuf_size2_399_out),
		.router_wrap_IVCH_0(mux_tree_tapbuf_size2_400_out),
		.router_wrap_IVCH_1(mux_tree_tapbuf_size2_401_out),
		.router_wrap_IVCH_2(mux_tree_tapbuf_size2_402_out),
		.router_wrap_IVCH_3(mux_tree_tapbuf_size2_403_out),
		.router_wrap_IVCH_4(mux_tree_tapbuf_size2_404_out),
		.router_wrap_IACK_0({mux_tree_tapbuf_size2_405_out, mux_tree_tapbuf_size2_406_out}),
		.router_wrap_IACK_1({mux_tree_tapbuf_size2_407_out, mux_tree_tapbuf_size2_408_out}),
		.router_wrap_IACK_2({mux_tree_tapbuf_size2_409_out, mux_tree_tapbuf_size2_410_out}),
		.router_wrap_IACK_3({mux_tree_tapbuf_size2_411_out, mux_tree_tapbuf_size2_412_out}),
		.router_wrap_IACK_4({mux_tree_tapbuf_size2_413_out, mux_tree_tapbuf_size2_414_out}),
		.router_wrap_ILCK_0({mux_tree_tapbuf_size2_415_out, mux_tree_tapbuf_size2_416_out}),
		.router_wrap_ILCK_1({mux_tree_tapbuf_size2_417_out, mux_tree_tapbuf_size2_418_out}),
		.router_wrap_ILCK_2({mux_tree_tapbuf_size2_419_out, mux_tree_tapbuf_size2_420_out}),
		.router_wrap_ILCK_3({mux_tree_tapbuf_size2_421_out, mux_tree_tapbuf_size2_422_out}),
		.router_wrap_ILCK_4({mux_tree_tapbuf_size2_423_out, mux_tree_tapbuf_size2_424_out}),
		.router_wrap_ODATA_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[0:34]),
		.router_wrap_ODATA_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[0:34]),
		.router_wrap_ODATA_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[0:34]),
		.router_wrap_ODATA_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[0:34]),
		.router_wrap_ODATA_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[0:34]),
		.router_wrap_OVALID_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_0),
		.router_wrap_OVALID_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_1),
		.router_wrap_OVALID_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_2),
		.router_wrap_OVALID_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_3),
		.router_wrap_OVALID_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_4),
		.router_wrap_OVCH_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_0),
		.router_wrap_OVCH_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_1),
		.router_wrap_OVCH_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_2),
		.router_wrap_OVCH_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_3),
		.router_wrap_OVCH_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_4),
		.router_wrap_OACK_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0[0:1]),
		.router_wrap_OACK_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1[0:1]),
		.router_wrap_OACK_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2[0:1]),
		.router_wrap_OACK_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3[0:1]),
		.router_wrap_OACK_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4[0:1]),
		.router_wrap_ORDY_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0[0:1]),
		.router_wrap_ORDY_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1[0:1]),
		.router_wrap_ORDY_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2[0:1]),
		.router_wrap_ORDY_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3[0:1]),
		.router_wrap_ORDY_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4[0:1]),
		.router_wrap_OLCK_0(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0[0:1]),
		.router_wrap_OLCK_1(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1[0:1]),
		.router_wrap_OLCK_2(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2[0:1]),
		.router_wrap_OLCK_3(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3[0:1]),
		.router_wrap_OLCK_4(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4[0:1]));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_RST_ logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_RST__0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_RST__D(direct_interc_0_out),
		.ff_RST__Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_RST__0_ff_RST__Q),
		.ff_RST__clk(direct_interc_1_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_MY_XPOS_D(direct_interc_2_out),
		.ff_MY_XPOS_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_0_ff_MY_XPOS_Q),
		.ff_MY_XPOS_clk(direct_interc_3_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_MY_XPOS_D(direct_interc_4_out),
		.ff_MY_XPOS_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_1_ff_MY_XPOS_Q),
		.ff_MY_XPOS_clk(direct_interc_5_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_MY_YPOS_D(direct_interc_6_out),
		.ff_MY_YPOS_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_0_ff_MY_YPOS_Q),
		.ff_MY_YPOS_clk(direct_interc_7_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_MY_YPOS_D(direct_interc_8_out),
		.ff_MY_YPOS_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_1_ff_MY_YPOS_Q),
		.ff_MY_YPOS_clk(direct_interc_9_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_10_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_0_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_11_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_12_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_1_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_13_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_14_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_2_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_15_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_16_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_3_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_17_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_18_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_4_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_19_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_20_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_5_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_21_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_22_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_6_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_23_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_24_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_7_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_25_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_26_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_8_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_27_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_28_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_9_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_29_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_30_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_10_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_31_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_32_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_11_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_33_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_34_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_12_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_35_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_36_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_13_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_37_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_38_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_14_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_39_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_40_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_15_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_41_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_42_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_16_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_43_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_44_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_17_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_45_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_46_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_18_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_47_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_48_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_19_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_49_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_50_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_20_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_51_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_52_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_21_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_53_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_54_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_22_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_55_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_56_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_23_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_57_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_58_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_24_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_59_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_60_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_25_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_61_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_62_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_26_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_63_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_64_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_27_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_65_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_66_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_28_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_67_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_68_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_29_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_69_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_70_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_30_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_71_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_72_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_31_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_73_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_74_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_32_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_75_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_76_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_33_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_77_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_0_D(direct_interc_78_out),
		.ff_IDATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_34_ff_IDATA_0_Q),
		.ff_IDATA_0_clk(direct_interc_79_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_80_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_0_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_81_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_82_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_1_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_83_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_84_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_2_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_85_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_86_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_3_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_87_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_88_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_4_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_89_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_90_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_5_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_91_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_92_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_6_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_93_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_94_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_7_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_95_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_96_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_8_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_97_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_98_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_9_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_99_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_100_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_10_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_101_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_102_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_11_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_103_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_104_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_12_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_105_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_106_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_13_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_107_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_108_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_14_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_109_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_110_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_15_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_111_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_112_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_16_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_113_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_114_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_17_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_115_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_116_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_18_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_117_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_118_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_19_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_119_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_120_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_20_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_121_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_122_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_21_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_123_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_124_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_22_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_125_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_126_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_23_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_127_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_128_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_24_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_129_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_130_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_25_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_131_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_132_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_26_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_133_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_134_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_27_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_135_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_136_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_28_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_137_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_138_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_29_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_139_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_140_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_30_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_141_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_142_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_31_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_143_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_144_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_32_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_145_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_146_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_33_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_147_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_1_D(direct_interc_148_out),
		.ff_IDATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_34_ff_IDATA_1_Q),
		.ff_IDATA_1_clk(direct_interc_149_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_150_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_0_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_151_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_152_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_1_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_153_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_154_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_2_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_155_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_156_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_3_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_157_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_158_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_4_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_159_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_160_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_5_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_161_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_162_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_6_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_163_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_164_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_7_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_165_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_166_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_8_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_167_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_168_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_9_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_169_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_170_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_10_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_171_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_172_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_11_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_173_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_174_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_12_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_175_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_176_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_13_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_177_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_178_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_14_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_179_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_180_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_15_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_181_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_182_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_16_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_183_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_184_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_17_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_185_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_186_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_18_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_187_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_188_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_19_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_189_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_190_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_20_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_191_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_192_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_21_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_193_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_194_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_22_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_195_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_196_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_23_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_197_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_198_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_24_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_199_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_200_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_25_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_201_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_202_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_26_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_203_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_204_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_27_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_205_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_206_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_28_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_207_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_208_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_29_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_209_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_210_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_30_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_211_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_212_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_31_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_213_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_214_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_32_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_215_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_216_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_33_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_217_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_2_D(direct_interc_218_out),
		.ff_IDATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_34_ff_IDATA_2_Q),
		.ff_IDATA_2_clk(direct_interc_219_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_220_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_0_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_221_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_222_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_1_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_223_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_224_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_2_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_225_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_226_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_3_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_227_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_228_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_4_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_229_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_230_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_5_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_231_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_232_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_6_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_233_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_234_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_7_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_235_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_236_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_8_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_237_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_238_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_9_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_239_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_240_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_10_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_241_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_242_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_11_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_243_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_244_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_12_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_245_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_246_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_13_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_247_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_248_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_14_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_249_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_250_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_15_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_251_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_252_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_16_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_253_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_254_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_17_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_255_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_256_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_18_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_257_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_258_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_19_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_259_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_260_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_20_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_261_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_262_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_21_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_263_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_264_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_22_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_265_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_266_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_23_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_267_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_268_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_24_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_269_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_270_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_25_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_271_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_272_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_26_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_273_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_274_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_27_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_275_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_276_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_28_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_277_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_278_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_29_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_279_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_280_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_30_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_281_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_282_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_31_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_283_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_284_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_32_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_285_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_286_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_33_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_287_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_3_D(direct_interc_288_out),
		.ff_IDATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_34_ff_IDATA_3_Q),
		.ff_IDATA_3_clk(direct_interc_289_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_290_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_0_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_291_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_292_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_1_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_293_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_294_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_2_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_295_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_296_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_3_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_297_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_298_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_4_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_299_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_300_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_5_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_301_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_302_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_6_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_303_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_304_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_7_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_305_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_306_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_8_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_307_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_308_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_9_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_309_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_310_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_10_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_311_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_312_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_11_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_313_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_314_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_12_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_315_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_316_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_13_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_317_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_318_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_14_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_319_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_320_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_15_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_321_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_322_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_16_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_323_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_324_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_17_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_325_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_326_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_18_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_327_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_328_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_19_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_329_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_330_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_20_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_331_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_332_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_21_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_333_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_334_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_22_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_335_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_336_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_23_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_337_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_338_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_24_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_339_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_340_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_25_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_341_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_342_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_26_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_343_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_344_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_27_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_345_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_346_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_28_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_347_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_348_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_29_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_349_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_350_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_30_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_351_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_352_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_31_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_353_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_354_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_32_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_355_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_356_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_33_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_357_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IDATA_4_D(direct_interc_358_out),
		.ff_IDATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_34_ff_IDATA_4_Q),
		.ff_IDATA_4_clk(direct_interc_359_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVALID_0_D(direct_interc_360_out),
		.ff_IVALID_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_0_0_ff_IVALID_0_Q),
		.ff_IVALID_0_clk(direct_interc_361_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVALID_1_D(direct_interc_362_out),
		.ff_IVALID_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_1_0_ff_IVALID_1_Q),
		.ff_IVALID_1_clk(direct_interc_363_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVALID_2_D(direct_interc_364_out),
		.ff_IVALID_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_2_0_ff_IVALID_2_Q),
		.ff_IVALID_2_clk(direct_interc_365_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVALID_3_D(direct_interc_366_out),
		.ff_IVALID_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_3_0_ff_IVALID_3_Q),
		.ff_IVALID_3_clk(direct_interc_367_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVALID_4_D(direct_interc_368_out),
		.ff_IVALID_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_4_0_ff_IVALID_4_Q),
		.ff_IVALID_4_clk(direct_interc_369_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVCH_0_D(direct_interc_370_out),
		.ff_IVCH_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_0_0_ff_IVCH_0_Q),
		.ff_IVCH_0_clk(direct_interc_371_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVCH_1_D(direct_interc_372_out),
		.ff_IVCH_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_1_0_ff_IVCH_1_Q),
		.ff_IVCH_1_clk(direct_interc_373_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVCH_2_D(direct_interc_374_out),
		.ff_IVCH_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_2_0_ff_IVCH_2_Q),
		.ff_IVCH_2_clk(direct_interc_375_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVCH_3_D(direct_interc_376_out),
		.ff_IVCH_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_3_0_ff_IVCH_3_Q),
		.ff_IVCH_3_clk(direct_interc_377_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IVCH_4_D(direct_interc_378_out),
		.ff_IVCH_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_4_0_ff_IVCH_4_Q),
		.ff_IVCH_4_clk(direct_interc_379_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_0_D(direct_interc_380_out),
		.ff_IACK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_0_ff_IACK_0_Q),
		.ff_IACK_0_clk(direct_interc_381_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_0_D(direct_interc_382_out),
		.ff_IACK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_1_ff_IACK_0_Q),
		.ff_IACK_0_clk(direct_interc_383_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_1_D(direct_interc_384_out),
		.ff_IACK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_0_ff_IACK_1_Q),
		.ff_IACK_1_clk(direct_interc_385_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_1_D(direct_interc_386_out),
		.ff_IACK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_1_ff_IACK_1_Q),
		.ff_IACK_1_clk(direct_interc_387_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_2_D(direct_interc_388_out),
		.ff_IACK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_0_ff_IACK_2_Q),
		.ff_IACK_2_clk(direct_interc_389_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_2_D(direct_interc_390_out),
		.ff_IACK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_1_ff_IACK_2_Q),
		.ff_IACK_2_clk(direct_interc_391_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_3_D(direct_interc_392_out),
		.ff_IACK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_0_ff_IACK_3_Q),
		.ff_IACK_3_clk(direct_interc_393_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_3_D(direct_interc_394_out),
		.ff_IACK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_1_ff_IACK_3_Q),
		.ff_IACK_3_clk(direct_interc_395_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_4_D(direct_interc_396_out),
		.ff_IACK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_0_ff_IACK_4_Q),
		.ff_IACK_4_clk(direct_interc_397_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_IACK_4_D(direct_interc_398_out),
		.ff_IACK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_1_ff_IACK_4_Q),
		.ff_IACK_4_clk(direct_interc_399_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_0_D(direct_interc_400_out),
		.ff_ILCK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_0_ff_ILCK_0_Q),
		.ff_ILCK_0_clk(direct_interc_401_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_0_D(direct_interc_402_out),
		.ff_ILCK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_1_ff_ILCK_0_Q),
		.ff_ILCK_0_clk(direct_interc_403_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_1_D(direct_interc_404_out),
		.ff_ILCK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_0_ff_ILCK_1_Q),
		.ff_ILCK_1_clk(direct_interc_405_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_1_D(direct_interc_406_out),
		.ff_ILCK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_1_ff_ILCK_1_Q),
		.ff_ILCK_1_clk(direct_interc_407_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_2_D(direct_interc_408_out),
		.ff_ILCK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_0_ff_ILCK_2_Q),
		.ff_ILCK_2_clk(direct_interc_409_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_2_D(direct_interc_410_out),
		.ff_ILCK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_1_ff_ILCK_2_Q),
		.ff_ILCK_2_clk(direct_interc_411_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_3_D(direct_interc_412_out),
		.ff_ILCK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_0_ff_ILCK_3_Q),
		.ff_ILCK_3_clk(direct_interc_413_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_3_D(direct_interc_414_out),
		.ff_ILCK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_1_ff_ILCK_3_Q),
		.ff_ILCK_3_clk(direct_interc_415_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_4_D(direct_interc_416_out),
		.ff_ILCK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_0_ff_ILCK_4_Q),
		.ff_ILCK_4_clk(direct_interc_417_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ILCK_4_D(direct_interc_418_out),
		.ff_ILCK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_1_ff_ILCK_4_Q),
		.ff_ILCK_4_clk(direct_interc_419_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_420_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_0_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_421_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_422_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_1_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_423_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_424_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_2_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_425_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_426_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_3_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_427_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_428_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_4_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_429_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_430_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_5_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_431_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_432_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_6_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_433_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_434_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_7_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_435_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_436_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_8_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_437_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_438_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_9_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_439_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_440_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_10_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_441_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_442_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_11_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_443_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_444_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_12_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_445_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_446_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_13_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_447_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_448_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_14_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_449_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_450_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_15_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_451_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_452_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_16_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_453_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_454_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_17_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_455_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_456_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_18_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_457_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_458_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_19_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_459_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_460_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_20_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_461_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_462_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_21_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_463_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_464_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_22_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_465_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_466_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_23_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_467_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_468_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_24_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_469_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_470_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_25_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_471_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_472_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_26_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_473_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_474_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_27_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_475_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_476_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_28_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_477_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_478_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_29_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_479_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_480_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_30_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_481_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_482_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_31_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_483_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_484_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_32_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_485_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_486_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_33_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_487_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_0_D(direct_interc_488_out),
		.ff_ODATA_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_34_ff_ODATA_0_Q),
		.ff_ODATA_0_clk(direct_interc_489_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_490_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_0_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_491_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_492_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_1_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_493_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_494_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_2_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_495_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_496_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_3_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_497_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_498_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_4_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_499_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_500_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_5_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_501_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_502_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_6_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_503_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_504_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_7_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_505_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_506_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_8_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_507_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_508_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_9_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_509_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_510_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_10_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_511_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_512_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_11_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_513_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_514_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_12_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_515_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_516_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_13_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_517_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_518_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_14_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_519_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_520_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_15_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_521_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_522_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_16_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_523_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_524_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_17_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_525_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_526_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_18_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_527_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_528_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_19_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_529_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_530_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_20_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_531_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_532_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_21_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_533_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_534_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_22_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_535_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_536_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_23_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_537_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_538_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_24_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_539_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_540_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_25_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_541_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_542_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_26_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_543_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_544_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_27_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_545_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_546_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_28_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_547_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_548_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_29_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_549_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_550_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_30_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_551_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_552_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_31_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_553_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_554_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_32_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_555_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_556_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_33_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_557_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_1_D(direct_interc_558_out),
		.ff_ODATA_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_34_ff_ODATA_1_Q),
		.ff_ODATA_1_clk(direct_interc_559_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_560_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_0_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_561_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_562_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_1_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_563_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_564_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_2_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_565_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_566_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_3_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_567_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_568_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_4_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_569_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_570_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_5_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_571_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_572_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_6_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_573_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_574_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_7_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_575_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_576_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_8_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_577_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_578_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_9_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_579_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_580_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_10_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_581_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_582_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_11_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_583_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_584_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_12_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_585_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_586_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_13_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_587_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_588_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_14_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_589_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_590_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_15_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_591_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_592_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_16_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_593_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_594_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_17_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_595_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_596_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_18_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_597_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_598_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_19_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_599_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_600_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_20_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_601_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_602_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_21_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_603_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_604_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_22_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_605_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_606_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_23_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_607_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_608_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_24_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_609_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_610_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_25_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_611_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_612_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_26_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_613_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_614_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_27_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_615_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_616_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_28_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_617_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_618_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_29_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_619_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_620_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_30_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_621_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_622_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_31_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_623_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_624_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_32_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_625_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_626_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_33_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_627_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_2_D(direct_interc_628_out),
		.ff_ODATA_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_34_ff_ODATA_2_Q),
		.ff_ODATA_2_clk(direct_interc_629_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_630_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_0_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_631_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_632_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_1_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_633_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_634_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_2_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_635_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_636_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_3_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_637_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_638_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_4_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_639_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_640_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_5_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_641_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_642_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_6_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_643_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_644_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_7_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_645_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_646_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_8_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_647_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_648_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_9_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_649_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_650_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_10_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_651_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_652_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_11_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_653_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_654_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_12_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_655_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_656_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_13_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_657_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_658_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_14_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_659_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_660_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_15_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_661_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_662_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_16_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_663_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_664_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_17_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_665_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_666_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_18_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_667_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_668_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_19_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_669_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_670_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_20_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_671_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_672_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_21_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_673_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_674_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_22_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_675_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_676_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_23_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_677_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_678_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_24_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_679_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_680_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_25_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_681_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_682_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_26_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_683_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_684_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_27_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_685_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_686_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_28_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_687_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_688_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_29_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_689_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_690_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_30_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_691_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_692_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_31_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_693_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_694_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_32_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_695_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_696_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_33_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_697_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_3_D(direct_interc_698_out),
		.ff_ODATA_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_34_ff_ODATA_3_Q),
		.ff_ODATA_3_clk(direct_interc_699_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_700_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_0_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_701_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_702_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_1_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_703_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_2 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_704_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_2_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_705_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_3 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_706_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_3_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_707_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_4 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_708_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_4_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_709_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_5 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_710_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_5_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_711_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_6 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_712_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_6_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_713_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_7 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_714_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_7_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_715_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_8 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_716_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_8_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_717_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_9 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_718_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_9_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_719_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_10 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_720_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_10_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_721_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_11 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_722_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_11_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_723_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_12 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_724_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_12_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_725_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_13 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_726_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_13_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_727_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_14 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_728_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_14_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_729_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_15 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_730_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_15_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_731_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_16 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_732_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_16_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_733_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_17 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_734_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_17_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_735_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_18 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_736_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_18_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_737_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_19 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_738_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_19_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_739_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_20 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_740_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_20_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_741_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_21 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_742_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_21_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_743_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_22 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_744_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_22_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_745_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_23 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_746_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_23_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_747_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_24 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_748_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_24_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_749_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_25 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_750_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_25_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_751_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_26 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_752_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_26_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_753_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_27 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_754_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_27_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_755_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_28 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_756_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_28_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_757_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_29 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_758_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_29_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_759_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_30 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_760_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_30_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_761_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_31 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_762_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_31_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_763_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_32 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_764_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_32_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_765_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_33 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_766_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_33_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_767_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_34 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ODATA_4_D(direct_interc_768_out),
		.ff_ODATA_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_34_ff_ODATA_4_Q),
		.ff_ODATA_4_clk(direct_interc_769_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVALID_0_D(direct_interc_770_out),
		.ff_OVALID_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_0_0_ff_OVALID_0_Q),
		.ff_OVALID_0_clk(direct_interc_771_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVALID_1_D(direct_interc_772_out),
		.ff_OVALID_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_1_0_ff_OVALID_1_Q),
		.ff_OVALID_1_clk(direct_interc_773_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVALID_2_D(direct_interc_774_out),
		.ff_OVALID_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_2_0_ff_OVALID_2_Q),
		.ff_OVALID_2_clk(direct_interc_775_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVALID_3_D(direct_interc_776_out),
		.ff_OVALID_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_3_0_ff_OVALID_3_Q),
		.ff_OVALID_3_clk(direct_interc_777_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVALID_4_D(direct_interc_778_out),
		.ff_OVALID_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_4_0_ff_OVALID_4_Q),
		.ff_OVALID_4_clk(direct_interc_779_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVCH_0_D(direct_interc_780_out),
		.ff_OVCH_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_0_0_ff_OVCH_0_Q),
		.ff_OVCH_0_clk(direct_interc_781_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVCH_1_D(direct_interc_782_out),
		.ff_OVCH_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_1_0_ff_OVCH_1_Q),
		.ff_OVCH_1_clk(direct_interc_783_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVCH_2_D(direct_interc_784_out),
		.ff_OVCH_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_2_0_ff_OVCH_2_Q),
		.ff_OVCH_2_clk(direct_interc_785_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVCH_3_D(direct_interc_786_out),
		.ff_OVCH_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_3_0_ff_OVCH_3_Q),
		.ff_OVCH_3_clk(direct_interc_787_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OVCH_4_D(direct_interc_788_out),
		.ff_OVCH_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_4_0_ff_OVCH_4_Q),
		.ff_OVCH_4_clk(direct_interc_789_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_0_D(direct_interc_790_out),
		.ff_OACK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_0_ff_OACK_0_Q),
		.ff_OACK_0_clk(direct_interc_791_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_0_D(direct_interc_792_out),
		.ff_OACK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_1_ff_OACK_0_Q),
		.ff_OACK_0_clk(direct_interc_793_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_1_D(direct_interc_794_out),
		.ff_OACK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_0_ff_OACK_1_Q),
		.ff_OACK_1_clk(direct_interc_795_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_1_D(direct_interc_796_out),
		.ff_OACK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_1_ff_OACK_1_Q),
		.ff_OACK_1_clk(direct_interc_797_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_2_D(direct_interc_798_out),
		.ff_OACK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_0_ff_OACK_2_Q),
		.ff_OACK_2_clk(direct_interc_799_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_2_D(direct_interc_800_out),
		.ff_OACK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_1_ff_OACK_2_Q),
		.ff_OACK_2_clk(direct_interc_801_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_3_D(direct_interc_802_out),
		.ff_OACK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_0_ff_OACK_3_Q),
		.ff_OACK_3_clk(direct_interc_803_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_3_D(direct_interc_804_out),
		.ff_OACK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_1_ff_OACK_3_Q),
		.ff_OACK_3_clk(direct_interc_805_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_4_D(direct_interc_806_out),
		.ff_OACK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_0_ff_OACK_4_Q),
		.ff_OACK_4_clk(direct_interc_807_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OACK_4_D(direct_interc_808_out),
		.ff_OACK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_1_ff_OACK_4_Q),
		.ff_OACK_4_clk(direct_interc_809_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_0_D(direct_interc_810_out),
		.ff_ORDY_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_0_ff_ORDY_0_Q),
		.ff_ORDY_0_clk(direct_interc_811_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_0_D(direct_interc_812_out),
		.ff_ORDY_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_1_ff_ORDY_0_Q),
		.ff_ORDY_0_clk(direct_interc_813_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_1_D(direct_interc_814_out),
		.ff_ORDY_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_0_ff_ORDY_1_Q),
		.ff_ORDY_1_clk(direct_interc_815_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_1_D(direct_interc_816_out),
		.ff_ORDY_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_1_ff_ORDY_1_Q),
		.ff_ORDY_1_clk(direct_interc_817_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_2_D(direct_interc_818_out),
		.ff_ORDY_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_0_ff_ORDY_2_Q),
		.ff_ORDY_2_clk(direct_interc_819_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_2_D(direct_interc_820_out),
		.ff_ORDY_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_1_ff_ORDY_2_Q),
		.ff_ORDY_2_clk(direct_interc_821_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_3_D(direct_interc_822_out),
		.ff_ORDY_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_0_ff_ORDY_3_Q),
		.ff_ORDY_3_clk(direct_interc_823_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_3_D(direct_interc_824_out),
		.ff_ORDY_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_1_ff_ORDY_3_Q),
		.ff_ORDY_3_clk(direct_interc_825_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_4_D(direct_interc_826_out),
		.ff_ORDY_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_0_ff_ORDY_4_Q),
		.ff_ORDY_4_clk(direct_interc_827_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_ORDY_4_D(direct_interc_828_out),
		.ff_ORDY_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_1_ff_ORDY_4_Q),
		.ff_ORDY_4_clk(direct_interc_829_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_0_D(direct_interc_830_out),
		.ff_OLCK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_0_ff_OLCK_0_Q),
		.ff_OLCK_0_clk(direct_interc_831_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_0_D(direct_interc_832_out),
		.ff_OLCK_0_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_1_ff_OLCK_0_Q),
		.ff_OLCK_0_clk(direct_interc_833_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_1_D(direct_interc_834_out),
		.ff_OLCK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_0_ff_OLCK_1_Q),
		.ff_OLCK_1_clk(direct_interc_835_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_1_D(direct_interc_836_out),
		.ff_OLCK_1_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_1_ff_OLCK_1_Q),
		.ff_OLCK_1_clk(direct_interc_837_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_2_D(direct_interc_838_out),
		.ff_OLCK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_0_ff_OLCK_2_Q),
		.ff_OLCK_2_clk(direct_interc_839_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_2_D(direct_interc_840_out),
		.ff_OLCK_2_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_1_ff_OLCK_2_Q),
		.ff_OLCK_2_clk(direct_interc_841_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_3_D(direct_interc_842_out),
		.ff_OLCK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_0_ff_OLCK_3_Q),
		.ff_OLCK_3_clk(direct_interc_843_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_3_D(direct_interc_844_out),
		.ff_OLCK_3_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_1_ff_OLCK_3_Q),
		.ff_OLCK_3_clk(direct_interc_845_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_0 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_4_D(direct_interc_846_out),
		.ff_OLCK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_0_ff_OLCK_4_Q),
		.ff_OLCK_4_clk(direct_interc_847_out));

	logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4 logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_1 (
		.set(set),
		.reset(reset),
		.clk(clk),
		.ff_OLCK_4_D(direct_interc_848_out),
		.ff_OLCK_4_Q(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_1_ff_OLCK_4_Q),
		.ff_OLCK_4_clk(direct_interc_849_out));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_0_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_1_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_2 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_2_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[2]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_3 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_3_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[3]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_4 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_4_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[4]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_5 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_5_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[5]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_6 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_6_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[6]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_7 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_7_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[7]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_8 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_8_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[8]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_9 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_9_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[9]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_10 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_10_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[10]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_11 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_11_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[11]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_12 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_12_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[12]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_13 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_13_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[13]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_14 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_14_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[14]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_15 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_15_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[15]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_16 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_16_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[16]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_17 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_17_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[17]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_18 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_18_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[18]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_19 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_19_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[19]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_20 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_20_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[20]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_21 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_21_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[21]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_22 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_22_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[22]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_23 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_23_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[23]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_24 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_24_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[24]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_25 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_25_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[25]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_26 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_26_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[26]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_27 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_27_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[27]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_28 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_28_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[28]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_29 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_29_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[29]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_30 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_30_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[30]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_31 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_31_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[31]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_32 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_32_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[32]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_33 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_33_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[33]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_0_cfg_34 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_0_34_ff_ODATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_0_cfg[34]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_0_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_1_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_2 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_2_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[2]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_3 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_3_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[3]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_4 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_4_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[4]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_5 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_5_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_40_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[5]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_6 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_6_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_41_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[6]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_7 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_7_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_42_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[7]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_8 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_8_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_43_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[8]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_9 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_9_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_44_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[9]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_10 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_10_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_45_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[10]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_11 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_11_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_46_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[11]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_12 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_12_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_47_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[12]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_13 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_13_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_48_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[13]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_14 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_14_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_49_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[14]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_15 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_15_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_50_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[15]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_16 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_16_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_51_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[16]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_17 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_17_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_52_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[17]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_18 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_18_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_53_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[18]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_19 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_19_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_54_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[19]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_20 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_20_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_55_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[20]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_21 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_21_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_56_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[21]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_22 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_22_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_57_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[22]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_23 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_23_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_58_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[23]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_24 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_24_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_59_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[24]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_25 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_25_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_60_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[25]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_26 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_26_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_61_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[26]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_27 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_27_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_62_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[27]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_28 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_28_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_63_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[28]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_29 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_29_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_64_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[29]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_30 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_30_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_65_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[30]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_31 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_31_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_66_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[31]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_32 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_32_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_67_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[32]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_33 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_33_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_68_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[33]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_1_cfg_34 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_1_34_ff_ODATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_69_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_1_cfg[34]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_0_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_70_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_1_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_71_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_2 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_2_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_72_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[2]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_3 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_3_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_73_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[3]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_4 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_4_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_74_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[4]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_5 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_5_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_75_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[5]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_6 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_6_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_76_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[6]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_7 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_7_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_77_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[7]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_8 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_8_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_78_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[8]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_9 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_9_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_79_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[9]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_10 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_10_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_80_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[10]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_11 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_11_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_81_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[11]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_12 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_12_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_82_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[12]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_13 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_13_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_83_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[13]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_14 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_14_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_84_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[14]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_15 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_15_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_85_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[15]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_16 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_16_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_86_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[16]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_17 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_17_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_87_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[17]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_18 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_18_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_88_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[18]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_19 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_19_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_89_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[19]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_20 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_20_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_90_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[20]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_21 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_21_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_91_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[21]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_22 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_22_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_92_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[22]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_23 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_23_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_93_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[23]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_24 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_24_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_94_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[24]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_25 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_25_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_95_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[25]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_26 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_26_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_96_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[26]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_27 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_27_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_97_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[27]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_28 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_28_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_98_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[28]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_29 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_29_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_99_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[29]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_30 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_30_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_100_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[30]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_31 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_31_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_101_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[31]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_32 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_32_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_102_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[32]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_33 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_33_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_103_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[33]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_2_cfg_34 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_2_34_ff_ODATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_104_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_2_cfg[34]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_0_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_105_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_1_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_106_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_2 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_2_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_107_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[2]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_3 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_3_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_108_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[3]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_4 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_4_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_109_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[4]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_5 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_5_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_110_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[5]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_6 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_6_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_111_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[6]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_7 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_7_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_112_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[7]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_8 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_8_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_113_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[8]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_9 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_9_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_114_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[9]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_10 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_10_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_115_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[10]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_11 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_11_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_116_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[11]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_12 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_12_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_117_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[12]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_13 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_13_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_118_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[13]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_14 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_14_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_119_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[14]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_15 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_15_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_120_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[15]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_16 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_16_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_121_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[16]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_17 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_17_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_122_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[17]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_18 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_18_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_123_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[18]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_19 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_19_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_124_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[19]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_20 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_20_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_125_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[20]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_21 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_21_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_126_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[21]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_22 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_22_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_127_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[22]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_23 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_23_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_128_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[23]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_24 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_24_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_129_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[24]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_25 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_25_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_130_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[25]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_26 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_26_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_131_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[26]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_27 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_27_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_132_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[27]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_28 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_28_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_133_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[28]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_29 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_29_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_134_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[29]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_30 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_30_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_135_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[30]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_31 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_31_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_136_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[31]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_32 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_32_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_137_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_137_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[32]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_33 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_33_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_138_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_138_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[33]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_3_cfg_34 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_3_34_ff_ODATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_139_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_139_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_3_cfg[34]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_0_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_140_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_140_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_1_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_141_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_141_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_2 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_2_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_142_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_142_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[2]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_3 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_3_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_143_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_143_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[3]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_4 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_4_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_144_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_144_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[4]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_5 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_5_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_145_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_145_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[5]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_6 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_6_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_146_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_146_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[6]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_7 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_7_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_147_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_147_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[7]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_8 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_8_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_148_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_148_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[8]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_9 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_9_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_149_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_149_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[9]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_10 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_10_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_150_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_150_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[10]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_11 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_11_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_151_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_151_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[11]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_12 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_12_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_152_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_152_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[12]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_13 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_13_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_153_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_153_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[13]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_14 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_14_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_154_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_154_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[14]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_15 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_15_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_155_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_155_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[15]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_16 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_16_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_156_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_156_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[16]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_17 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_17_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_157_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_157_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[17]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_18 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_18_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_158_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_158_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[18]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_19 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_19_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_159_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_159_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[19]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_20 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_20_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_160_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_160_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[20]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_21 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_21_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_161_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_161_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[21]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_22 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_22_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_162_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_162_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[22]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_23 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_23_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_163_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_163_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[23]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_24 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_24_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_164_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_164_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[24]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_25 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_25_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_165_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_165_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[25]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_26 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_26_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_166_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_166_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[26]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_27 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_27_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_167_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_167_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[27]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_28 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_28_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_168_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_168_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[28]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_29 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_29_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_169_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_169_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[29]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_30 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_30_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_170_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_170_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[30]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_31 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_31_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_171_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_171_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[31]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_32 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_32_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_172_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_172_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[32]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_33 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_33_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_173_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_173_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[33]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ODATA_4_cfg_34 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ODATA_4_34_ff_ODATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_174_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_174_sram_inv[0:1]),
		.out(router_wrap_slice_ODATA_4_cfg[34]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVALID_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_0, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_0_0_ff_OVALID_0_Q}),
		.sram(mux_tree_tapbuf_size2_175_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_175_sram_inv[0:1]),
		.out(router_wrap_slice_OVALID_0_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVALID_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_1, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_1_0_ff_OVALID_1_Q}),
		.sram(mux_tree_tapbuf_size2_176_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_176_sram_inv[0:1]),
		.out(router_wrap_slice_OVALID_1_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVALID_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_2, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_2_0_ff_OVALID_2_Q}),
		.sram(mux_tree_tapbuf_size2_177_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_177_sram_inv[0:1]),
		.out(router_wrap_slice_OVALID_2_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVALID_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_3, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_3_0_ff_OVALID_3_Q}),
		.sram(mux_tree_tapbuf_size2_178_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_178_sram_inv[0:1]),
		.out(router_wrap_slice_OVALID_3_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVALID_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_4, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVALID_4_0_ff_OVALID_4_Q}),
		.sram(mux_tree_tapbuf_size2_179_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_179_sram_inv[0:1]),
		.out(router_wrap_slice_OVALID_4_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVCH_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_0, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_0_0_ff_OVCH_0_Q}),
		.sram(mux_tree_tapbuf_size2_180_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_180_sram_inv[0:1]),
		.out(router_wrap_slice_OVCH_0_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVCH_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_1, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_1_0_ff_OVCH_1_Q}),
		.sram(mux_tree_tapbuf_size2_181_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_181_sram_inv[0:1]),
		.out(router_wrap_slice_OVCH_1_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVCH_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_2, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_2_0_ff_OVCH_2_Q}),
		.sram(mux_tree_tapbuf_size2_182_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_182_sram_inv[0:1]),
		.out(router_wrap_slice_OVCH_2_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVCH_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_3, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_3_0_ff_OVCH_3_Q}),
		.sram(mux_tree_tapbuf_size2_183_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_183_sram_inv[0:1]),
		.out(router_wrap_slice_OVCH_3_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OVCH_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_4, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OVCH_4_0_ff_OVCH_4_Q}),
		.sram(mux_tree_tapbuf_size2_184_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_184_sram_inv[0:1]),
		.out(router_wrap_slice_OVCH_4_cfg));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_0_ff_OACK_0_Q}),
		.sram(mux_tree_tapbuf_size2_185_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_185_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_0_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_0_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_0_1_ff_OACK_0_Q}),
		.sram(mux_tree_tapbuf_size2_186_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_186_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_0_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_0_ff_OACK_1_Q}),
		.sram(mux_tree_tapbuf_size2_187_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_187_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_1_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_1_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_1_1_ff_OACK_1_Q}),
		.sram(mux_tree_tapbuf_size2_188_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_188_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_1_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_0_ff_OACK_2_Q}),
		.sram(mux_tree_tapbuf_size2_189_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_189_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_2_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_2_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_2_1_ff_OACK_2_Q}),
		.sram(mux_tree_tapbuf_size2_190_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_190_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_2_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_0_ff_OACK_3_Q}),
		.sram(mux_tree_tapbuf_size2_191_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_191_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_3_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_3_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_3_1_ff_OACK_3_Q}),
		.sram(mux_tree_tapbuf_size2_192_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_192_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_3_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_0_ff_OACK_4_Q}),
		.sram(mux_tree_tapbuf_size2_193_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_193_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_4_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OACK_4_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OACK_4_1_ff_OACK_4_Q}),
		.sram(mux_tree_tapbuf_size2_194_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_194_sram_inv[0:1]),
		.out(router_wrap_slice_OACK_4_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_0_ff_ORDY_0_Q}),
		.sram(mux_tree_tapbuf_size2_195_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_195_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_0_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_0_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_0_1_ff_ORDY_0_Q}),
		.sram(mux_tree_tapbuf_size2_196_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_196_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_0_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_0_ff_ORDY_1_Q}),
		.sram(mux_tree_tapbuf_size2_197_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_197_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_1_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_1_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_1_1_ff_ORDY_1_Q}),
		.sram(mux_tree_tapbuf_size2_198_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_198_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_1_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_0_ff_ORDY_2_Q}),
		.sram(mux_tree_tapbuf_size2_199_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_199_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_2_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_2_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_2_1_ff_ORDY_2_Q}),
		.sram(mux_tree_tapbuf_size2_200_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_200_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_2_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_0_ff_ORDY_3_Q}),
		.sram(mux_tree_tapbuf_size2_201_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_201_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_3_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_3_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_3_1_ff_ORDY_3_Q}),
		.sram(mux_tree_tapbuf_size2_202_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_202_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_3_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_0_ff_ORDY_4_Q}),
		.sram(mux_tree_tapbuf_size2_203_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_203_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_4_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_ORDY_4_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ORDY_4_1_ff_ORDY_4_Q}),
		.sram(mux_tree_tapbuf_size2_204_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_204_sram_inv[0:1]),
		.out(router_wrap_slice_ORDY_4_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_0_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_0_ff_OLCK_0_Q}),
		.sram(mux_tree_tapbuf_size2_205_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_205_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_0_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_0_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_0_1_ff_OLCK_0_Q}),
		.sram(mux_tree_tapbuf_size2_206_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_206_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_0_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_1_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_0_ff_OLCK_1_Q}),
		.sram(mux_tree_tapbuf_size2_207_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_207_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_1_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_1_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_1_1_ff_OLCK_1_Q}),
		.sram(mux_tree_tapbuf_size2_208_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_208_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_1_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_2_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_0_ff_OLCK_2_Q}),
		.sram(mux_tree_tapbuf_size2_209_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_209_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_2_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_2_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_2_1_ff_OLCK_2_Q}),
		.sram(mux_tree_tapbuf_size2_210_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_210_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_2_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_3_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_0_ff_OLCK_3_Q}),
		.sram(mux_tree_tapbuf_size2_211_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_211_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_3_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_3_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_3_1_ff_OLCK_3_Q}),
		.sram(mux_tree_tapbuf_size2_212_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_212_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_3_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_4_cfg_0 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_0_ff_OLCK_4_Q}),
		.sram(mux_tree_tapbuf_size2_213_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_213_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_4_cfg[0]));

	mux_tree_tapbuf_size2 mux_router_wrap_slice_OLCK_4_cfg_1 (
		.in({logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_OLCK_4_1_ff_OLCK_4_Q}),
		.sram(mux_tree_tapbuf_size2_214_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_214_sram_inv[0:1]),
		.out(router_wrap_slice_OLCK_4_cfg[1]));

	mux_tree_tapbuf_size2 mux_router_wrap_0_RST__0 (
		.in({router_wrap_slice_RST__cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_RST__0_ff_RST__Q}),
		.sram(mux_tree_tapbuf_size2_215_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_215_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_215_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_MY_XPOS_0 (
		.in({router_wrap_slice_MY_XPOS_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_0_ff_MY_XPOS_Q}),
		.sram(mux_tree_tapbuf_size2_216_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_216_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_216_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_MY_XPOS_1 (
		.in({router_wrap_slice_MY_XPOS_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_XPOS_1_ff_MY_XPOS_Q}),
		.sram(mux_tree_tapbuf_size2_217_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_217_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_217_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_MY_YPOS_0 (
		.in({router_wrap_slice_MY_YPOS_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_0_ff_MY_YPOS_Q}),
		.sram(mux_tree_tapbuf_size2_218_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_218_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_218_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_MY_YPOS_1 (
		.in({router_wrap_slice_MY_YPOS_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_MY_YPOS_1_ff_MY_YPOS_Q}),
		.sram(mux_tree_tapbuf_size2_219_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_219_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_219_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_0 (
		.in({router_wrap_slice_IDATA_0_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_0_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_220_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_220_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_220_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_1 (
		.in({router_wrap_slice_IDATA_0_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_1_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_221_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_221_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_221_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_2 (
		.in({router_wrap_slice_IDATA_0_cfg[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_2_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_222_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_222_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_222_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_3 (
		.in({router_wrap_slice_IDATA_0_cfg[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_3_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_223_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_223_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_223_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_4 (
		.in({router_wrap_slice_IDATA_0_cfg[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_4_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_224_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_224_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_224_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_5 (
		.in({router_wrap_slice_IDATA_0_cfg[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_5_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_225_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_225_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_225_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_6 (
		.in({router_wrap_slice_IDATA_0_cfg[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_6_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_226_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_226_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_226_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_7 (
		.in({router_wrap_slice_IDATA_0_cfg[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_7_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_227_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_227_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_227_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_8 (
		.in({router_wrap_slice_IDATA_0_cfg[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_8_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_228_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_228_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_228_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_9 (
		.in({router_wrap_slice_IDATA_0_cfg[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_9_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_229_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_229_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_229_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_10 (
		.in({router_wrap_slice_IDATA_0_cfg[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_10_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_230_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_230_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_230_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_11 (
		.in({router_wrap_slice_IDATA_0_cfg[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_11_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_231_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_231_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_231_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_12 (
		.in({router_wrap_slice_IDATA_0_cfg[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_12_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_232_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_232_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_232_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_13 (
		.in({router_wrap_slice_IDATA_0_cfg[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_13_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_233_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_233_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_233_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_14 (
		.in({router_wrap_slice_IDATA_0_cfg[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_14_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_234_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_234_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_234_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_15 (
		.in({router_wrap_slice_IDATA_0_cfg[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_15_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_235_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_235_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_235_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_16 (
		.in({router_wrap_slice_IDATA_0_cfg[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_16_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_236_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_236_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_236_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_17 (
		.in({router_wrap_slice_IDATA_0_cfg[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_17_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_237_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_237_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_237_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_18 (
		.in({router_wrap_slice_IDATA_0_cfg[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_18_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_238_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_238_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_238_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_19 (
		.in({router_wrap_slice_IDATA_0_cfg[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_19_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_239_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_239_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_239_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_20 (
		.in({router_wrap_slice_IDATA_0_cfg[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_20_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_240_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_240_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_240_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_21 (
		.in({router_wrap_slice_IDATA_0_cfg[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_21_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_241_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_241_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_241_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_22 (
		.in({router_wrap_slice_IDATA_0_cfg[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_22_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_242_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_242_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_242_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_23 (
		.in({router_wrap_slice_IDATA_0_cfg[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_23_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_243_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_243_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_243_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_24 (
		.in({router_wrap_slice_IDATA_0_cfg[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_24_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_244_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_244_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_244_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_25 (
		.in({router_wrap_slice_IDATA_0_cfg[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_25_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_245_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_245_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_245_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_26 (
		.in({router_wrap_slice_IDATA_0_cfg[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_26_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_246_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_246_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_246_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_27 (
		.in({router_wrap_slice_IDATA_0_cfg[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_27_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_247_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_247_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_247_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_28 (
		.in({router_wrap_slice_IDATA_0_cfg[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_28_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_248_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_248_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_248_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_29 (
		.in({router_wrap_slice_IDATA_0_cfg[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_29_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_249_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_249_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_249_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_30 (
		.in({router_wrap_slice_IDATA_0_cfg[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_30_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_250_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_250_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_250_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_31 (
		.in({router_wrap_slice_IDATA_0_cfg[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_31_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_251_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_251_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_251_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_32 (
		.in({router_wrap_slice_IDATA_0_cfg[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_32_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_252_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_252_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_252_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_33 (
		.in({router_wrap_slice_IDATA_0_cfg[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_33_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_253_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_253_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_253_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_0_34 (
		.in({router_wrap_slice_IDATA_0_cfg[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_0_34_ff_IDATA_0_Q}),
		.sram(mux_tree_tapbuf_size2_254_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_254_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_254_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_0 (
		.in({router_wrap_slice_IDATA_1_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_0_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_255_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_255_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_255_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_1 (
		.in({router_wrap_slice_IDATA_1_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_1_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_256_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_256_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_256_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_2 (
		.in({router_wrap_slice_IDATA_1_cfg[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_2_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_257_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_257_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_257_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_3 (
		.in({router_wrap_slice_IDATA_1_cfg[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_3_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_258_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_258_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_258_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_4 (
		.in({router_wrap_slice_IDATA_1_cfg[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_4_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_259_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_259_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_259_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_5 (
		.in({router_wrap_slice_IDATA_1_cfg[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_5_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_260_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_260_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_260_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_6 (
		.in({router_wrap_slice_IDATA_1_cfg[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_6_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_261_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_261_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_261_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_7 (
		.in({router_wrap_slice_IDATA_1_cfg[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_7_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_262_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_262_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_262_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_8 (
		.in({router_wrap_slice_IDATA_1_cfg[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_8_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_263_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_263_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_263_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_9 (
		.in({router_wrap_slice_IDATA_1_cfg[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_9_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_264_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_264_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_264_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_10 (
		.in({router_wrap_slice_IDATA_1_cfg[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_10_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_265_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_265_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_265_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_11 (
		.in({router_wrap_slice_IDATA_1_cfg[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_11_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_266_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_266_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_266_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_12 (
		.in({router_wrap_slice_IDATA_1_cfg[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_12_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_267_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_267_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_267_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_13 (
		.in({router_wrap_slice_IDATA_1_cfg[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_13_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_268_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_268_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_268_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_14 (
		.in({router_wrap_slice_IDATA_1_cfg[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_14_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_269_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_269_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_269_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_15 (
		.in({router_wrap_slice_IDATA_1_cfg[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_15_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_270_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_270_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_270_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_16 (
		.in({router_wrap_slice_IDATA_1_cfg[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_16_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_271_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_271_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_271_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_17 (
		.in({router_wrap_slice_IDATA_1_cfg[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_17_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_272_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_272_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_272_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_18 (
		.in({router_wrap_slice_IDATA_1_cfg[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_18_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_273_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_273_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_273_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_19 (
		.in({router_wrap_slice_IDATA_1_cfg[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_19_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_274_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_274_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_274_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_20 (
		.in({router_wrap_slice_IDATA_1_cfg[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_20_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_275_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_275_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_275_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_21 (
		.in({router_wrap_slice_IDATA_1_cfg[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_21_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_276_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_276_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_276_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_22 (
		.in({router_wrap_slice_IDATA_1_cfg[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_22_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_277_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_277_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_277_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_23 (
		.in({router_wrap_slice_IDATA_1_cfg[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_23_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_278_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_278_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_278_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_24 (
		.in({router_wrap_slice_IDATA_1_cfg[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_24_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_279_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_279_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_279_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_25 (
		.in({router_wrap_slice_IDATA_1_cfg[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_25_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_280_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_280_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_280_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_26 (
		.in({router_wrap_slice_IDATA_1_cfg[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_26_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_281_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_281_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_281_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_27 (
		.in({router_wrap_slice_IDATA_1_cfg[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_27_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_282_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_282_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_282_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_28 (
		.in({router_wrap_slice_IDATA_1_cfg[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_28_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_283_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_283_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_283_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_29 (
		.in({router_wrap_slice_IDATA_1_cfg[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_29_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_284_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_284_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_284_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_30 (
		.in({router_wrap_slice_IDATA_1_cfg[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_30_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_285_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_285_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_285_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_31 (
		.in({router_wrap_slice_IDATA_1_cfg[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_31_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_286_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_286_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_286_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_32 (
		.in({router_wrap_slice_IDATA_1_cfg[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_32_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_287_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_287_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_287_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_33 (
		.in({router_wrap_slice_IDATA_1_cfg[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_33_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_288_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_288_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_288_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_1_34 (
		.in({router_wrap_slice_IDATA_1_cfg[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_1_34_ff_IDATA_1_Q}),
		.sram(mux_tree_tapbuf_size2_289_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_289_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_289_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_0 (
		.in({router_wrap_slice_IDATA_2_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_0_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_290_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_290_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_290_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_1 (
		.in({router_wrap_slice_IDATA_2_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_1_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_291_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_291_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_291_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_2 (
		.in({router_wrap_slice_IDATA_2_cfg[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_2_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_292_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_292_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_292_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_3 (
		.in({router_wrap_slice_IDATA_2_cfg[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_3_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_293_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_293_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_293_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_4 (
		.in({router_wrap_slice_IDATA_2_cfg[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_4_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_294_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_294_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_294_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_5 (
		.in({router_wrap_slice_IDATA_2_cfg[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_5_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_295_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_295_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_295_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_6 (
		.in({router_wrap_slice_IDATA_2_cfg[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_6_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_296_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_296_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_296_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_7 (
		.in({router_wrap_slice_IDATA_2_cfg[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_7_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_297_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_297_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_297_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_8 (
		.in({router_wrap_slice_IDATA_2_cfg[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_8_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_298_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_298_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_298_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_9 (
		.in({router_wrap_slice_IDATA_2_cfg[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_9_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_299_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_299_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_299_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_10 (
		.in({router_wrap_slice_IDATA_2_cfg[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_10_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_300_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_300_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_300_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_11 (
		.in({router_wrap_slice_IDATA_2_cfg[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_11_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_301_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_301_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_301_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_12 (
		.in({router_wrap_slice_IDATA_2_cfg[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_12_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_302_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_302_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_302_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_13 (
		.in({router_wrap_slice_IDATA_2_cfg[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_13_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_303_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_303_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_303_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_14 (
		.in({router_wrap_slice_IDATA_2_cfg[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_14_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_304_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_304_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_304_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_15 (
		.in({router_wrap_slice_IDATA_2_cfg[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_15_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_305_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_305_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_305_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_16 (
		.in({router_wrap_slice_IDATA_2_cfg[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_16_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_306_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_306_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_306_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_17 (
		.in({router_wrap_slice_IDATA_2_cfg[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_17_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_307_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_307_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_307_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_18 (
		.in({router_wrap_slice_IDATA_2_cfg[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_18_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_308_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_308_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_308_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_19 (
		.in({router_wrap_slice_IDATA_2_cfg[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_19_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_309_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_309_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_309_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_20 (
		.in({router_wrap_slice_IDATA_2_cfg[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_20_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_310_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_310_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_310_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_21 (
		.in({router_wrap_slice_IDATA_2_cfg[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_21_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_311_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_311_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_311_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_22 (
		.in({router_wrap_slice_IDATA_2_cfg[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_22_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_312_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_312_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_312_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_23 (
		.in({router_wrap_slice_IDATA_2_cfg[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_23_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_313_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_313_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_313_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_24 (
		.in({router_wrap_slice_IDATA_2_cfg[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_24_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_314_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_314_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_314_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_25 (
		.in({router_wrap_slice_IDATA_2_cfg[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_25_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_315_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_315_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_315_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_26 (
		.in({router_wrap_slice_IDATA_2_cfg[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_26_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_316_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_316_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_316_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_27 (
		.in({router_wrap_slice_IDATA_2_cfg[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_27_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_317_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_317_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_317_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_28 (
		.in({router_wrap_slice_IDATA_2_cfg[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_28_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_318_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_318_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_318_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_29 (
		.in({router_wrap_slice_IDATA_2_cfg[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_29_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_319_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_319_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_319_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_30 (
		.in({router_wrap_slice_IDATA_2_cfg[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_30_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_320_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_320_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_320_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_31 (
		.in({router_wrap_slice_IDATA_2_cfg[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_31_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_321_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_321_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_321_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_32 (
		.in({router_wrap_slice_IDATA_2_cfg[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_32_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_322_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_322_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_322_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_33 (
		.in({router_wrap_slice_IDATA_2_cfg[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_33_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_323_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_323_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_323_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_2_34 (
		.in({router_wrap_slice_IDATA_2_cfg[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_2_34_ff_IDATA_2_Q}),
		.sram(mux_tree_tapbuf_size2_324_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_324_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_324_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_0 (
		.in({router_wrap_slice_IDATA_3_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_0_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_325_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_325_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_325_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_1 (
		.in({router_wrap_slice_IDATA_3_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_1_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_326_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_326_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_326_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_2 (
		.in({router_wrap_slice_IDATA_3_cfg[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_2_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_327_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_327_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_327_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_3 (
		.in({router_wrap_slice_IDATA_3_cfg[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_3_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_328_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_328_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_328_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_4 (
		.in({router_wrap_slice_IDATA_3_cfg[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_4_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_329_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_329_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_329_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_5 (
		.in({router_wrap_slice_IDATA_3_cfg[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_5_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_330_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_330_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_330_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_6 (
		.in({router_wrap_slice_IDATA_3_cfg[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_6_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_331_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_331_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_331_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_7 (
		.in({router_wrap_slice_IDATA_3_cfg[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_7_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_332_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_332_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_332_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_8 (
		.in({router_wrap_slice_IDATA_3_cfg[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_8_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_333_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_333_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_333_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_9 (
		.in({router_wrap_slice_IDATA_3_cfg[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_9_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_334_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_334_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_334_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_10 (
		.in({router_wrap_slice_IDATA_3_cfg[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_10_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_335_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_335_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_335_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_11 (
		.in({router_wrap_slice_IDATA_3_cfg[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_11_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_336_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_336_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_336_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_12 (
		.in({router_wrap_slice_IDATA_3_cfg[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_12_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_337_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_337_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_337_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_13 (
		.in({router_wrap_slice_IDATA_3_cfg[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_13_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_338_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_338_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_338_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_14 (
		.in({router_wrap_slice_IDATA_3_cfg[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_14_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_339_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_339_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_339_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_15 (
		.in({router_wrap_slice_IDATA_3_cfg[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_15_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_340_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_340_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_340_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_16 (
		.in({router_wrap_slice_IDATA_3_cfg[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_16_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_341_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_341_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_341_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_17 (
		.in({router_wrap_slice_IDATA_3_cfg[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_17_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_342_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_342_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_342_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_18 (
		.in({router_wrap_slice_IDATA_3_cfg[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_18_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_343_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_343_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_343_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_19 (
		.in({router_wrap_slice_IDATA_3_cfg[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_19_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_344_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_344_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_344_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_20 (
		.in({router_wrap_slice_IDATA_3_cfg[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_20_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_345_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_345_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_345_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_21 (
		.in({router_wrap_slice_IDATA_3_cfg[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_21_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_346_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_346_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_346_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_22 (
		.in({router_wrap_slice_IDATA_3_cfg[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_22_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_347_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_347_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_347_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_23 (
		.in({router_wrap_slice_IDATA_3_cfg[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_23_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_348_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_348_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_348_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_24 (
		.in({router_wrap_slice_IDATA_3_cfg[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_24_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_349_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_349_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_349_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_25 (
		.in({router_wrap_slice_IDATA_3_cfg[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_25_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_350_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_350_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_350_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_26 (
		.in({router_wrap_slice_IDATA_3_cfg[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_26_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_351_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_351_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_351_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_27 (
		.in({router_wrap_slice_IDATA_3_cfg[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_27_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_352_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_352_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_352_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_28 (
		.in({router_wrap_slice_IDATA_3_cfg[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_28_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_353_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_353_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_353_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_29 (
		.in({router_wrap_slice_IDATA_3_cfg[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_29_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_354_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_354_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_354_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_30 (
		.in({router_wrap_slice_IDATA_3_cfg[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_30_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_355_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_355_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_355_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_31 (
		.in({router_wrap_slice_IDATA_3_cfg[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_31_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_356_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_356_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_356_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_32 (
		.in({router_wrap_slice_IDATA_3_cfg[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_32_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_357_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_357_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_357_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_33 (
		.in({router_wrap_slice_IDATA_3_cfg[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_33_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_358_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_358_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_358_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_3_34 (
		.in({router_wrap_slice_IDATA_3_cfg[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_3_34_ff_IDATA_3_Q}),
		.sram(mux_tree_tapbuf_size2_359_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_359_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_359_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_0 (
		.in({router_wrap_slice_IDATA_4_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_0_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_360_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_360_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_360_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_1 (
		.in({router_wrap_slice_IDATA_4_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_1_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_361_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_361_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_361_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_2 (
		.in({router_wrap_slice_IDATA_4_cfg[2], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_2_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_362_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_362_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_362_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_3 (
		.in({router_wrap_slice_IDATA_4_cfg[3], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_3_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_363_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_363_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_363_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_4 (
		.in({router_wrap_slice_IDATA_4_cfg[4], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_4_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_364_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_364_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_364_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_5 (
		.in({router_wrap_slice_IDATA_4_cfg[5], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_5_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_365_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_365_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_365_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_6 (
		.in({router_wrap_slice_IDATA_4_cfg[6], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_6_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_366_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_366_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_366_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_7 (
		.in({router_wrap_slice_IDATA_4_cfg[7], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_7_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_367_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_367_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_367_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_8 (
		.in({router_wrap_slice_IDATA_4_cfg[8], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_8_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_368_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_368_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_368_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_9 (
		.in({router_wrap_slice_IDATA_4_cfg[9], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_9_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_369_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_369_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_369_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_10 (
		.in({router_wrap_slice_IDATA_4_cfg[10], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_10_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_370_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_370_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_370_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_11 (
		.in({router_wrap_slice_IDATA_4_cfg[11], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_11_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_371_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_371_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_371_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_12 (
		.in({router_wrap_slice_IDATA_4_cfg[12], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_12_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_372_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_372_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_372_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_13 (
		.in({router_wrap_slice_IDATA_4_cfg[13], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_13_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_373_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_373_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_373_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_14 (
		.in({router_wrap_slice_IDATA_4_cfg[14], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_14_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_374_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_374_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_374_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_15 (
		.in({router_wrap_slice_IDATA_4_cfg[15], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_15_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_375_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_375_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_375_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_16 (
		.in({router_wrap_slice_IDATA_4_cfg[16], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_16_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_376_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_376_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_376_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_17 (
		.in({router_wrap_slice_IDATA_4_cfg[17], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_17_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_377_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_377_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_377_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_18 (
		.in({router_wrap_slice_IDATA_4_cfg[18], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_18_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_378_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_378_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_378_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_19 (
		.in({router_wrap_slice_IDATA_4_cfg[19], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_19_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_379_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_379_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_379_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_20 (
		.in({router_wrap_slice_IDATA_4_cfg[20], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_20_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_380_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_380_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_380_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_21 (
		.in({router_wrap_slice_IDATA_4_cfg[21], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_21_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_381_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_381_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_381_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_22 (
		.in({router_wrap_slice_IDATA_4_cfg[22], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_22_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_382_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_382_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_382_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_23 (
		.in({router_wrap_slice_IDATA_4_cfg[23], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_23_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_383_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_383_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_383_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_24 (
		.in({router_wrap_slice_IDATA_4_cfg[24], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_24_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_384_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_384_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_384_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_25 (
		.in({router_wrap_slice_IDATA_4_cfg[25], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_25_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_385_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_385_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_385_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_26 (
		.in({router_wrap_slice_IDATA_4_cfg[26], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_26_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_386_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_386_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_386_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_27 (
		.in({router_wrap_slice_IDATA_4_cfg[27], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_27_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_387_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_387_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_387_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_28 (
		.in({router_wrap_slice_IDATA_4_cfg[28], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_28_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_388_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_388_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_388_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_29 (
		.in({router_wrap_slice_IDATA_4_cfg[29], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_29_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_389_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_389_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_389_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_30 (
		.in({router_wrap_slice_IDATA_4_cfg[30], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_30_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_390_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_390_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_390_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_31 (
		.in({router_wrap_slice_IDATA_4_cfg[31], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_31_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_391_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_391_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_391_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_32 (
		.in({router_wrap_slice_IDATA_4_cfg[32], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_32_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_392_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_392_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_392_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_33 (
		.in({router_wrap_slice_IDATA_4_cfg[33], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_33_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_393_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_393_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_393_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IDATA_4_34 (
		.in({router_wrap_slice_IDATA_4_cfg[34], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IDATA_4_34_ff_IDATA_4_Q}),
		.sram(mux_tree_tapbuf_size2_394_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_394_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_394_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVALID_0_0 (
		.in({router_wrap_slice_IVALID_0_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_0_0_ff_IVALID_0_Q}),
		.sram(mux_tree_tapbuf_size2_395_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_395_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_395_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVALID_1_0 (
		.in({router_wrap_slice_IVALID_1_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_1_0_ff_IVALID_1_Q}),
		.sram(mux_tree_tapbuf_size2_396_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_396_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_396_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVALID_2_0 (
		.in({router_wrap_slice_IVALID_2_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_2_0_ff_IVALID_2_Q}),
		.sram(mux_tree_tapbuf_size2_397_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_397_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_397_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVALID_3_0 (
		.in({router_wrap_slice_IVALID_3_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_3_0_ff_IVALID_3_Q}),
		.sram(mux_tree_tapbuf_size2_398_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_398_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_398_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVALID_4_0 (
		.in({router_wrap_slice_IVALID_4_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVALID_4_0_ff_IVALID_4_Q}),
		.sram(mux_tree_tapbuf_size2_399_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_399_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_399_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVCH_0_0 (
		.in({router_wrap_slice_IVCH_0_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_0_0_ff_IVCH_0_Q}),
		.sram(mux_tree_tapbuf_size2_400_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_400_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_400_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVCH_1_0 (
		.in({router_wrap_slice_IVCH_1_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_1_0_ff_IVCH_1_Q}),
		.sram(mux_tree_tapbuf_size2_401_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_401_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_401_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVCH_2_0 (
		.in({router_wrap_slice_IVCH_2_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_2_0_ff_IVCH_2_Q}),
		.sram(mux_tree_tapbuf_size2_402_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_402_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_402_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVCH_3_0 (
		.in({router_wrap_slice_IVCH_3_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_3_0_ff_IVCH_3_Q}),
		.sram(mux_tree_tapbuf_size2_403_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_403_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_403_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IVCH_4_0 (
		.in({router_wrap_slice_IVCH_4_cfg, logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IVCH_4_0_ff_IVCH_4_Q}),
		.sram(mux_tree_tapbuf_size2_404_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_404_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_404_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_0_0 (
		.in({router_wrap_slice_IACK_0_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_0_ff_IACK_0_Q}),
		.sram(mux_tree_tapbuf_size2_405_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_405_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_405_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_0_1 (
		.in({router_wrap_slice_IACK_0_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_0_1_ff_IACK_0_Q}),
		.sram(mux_tree_tapbuf_size2_406_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_406_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_406_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_1_0 (
		.in({router_wrap_slice_IACK_1_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_0_ff_IACK_1_Q}),
		.sram(mux_tree_tapbuf_size2_407_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_407_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_407_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_1_1 (
		.in({router_wrap_slice_IACK_1_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_1_1_ff_IACK_1_Q}),
		.sram(mux_tree_tapbuf_size2_408_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_408_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_408_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_2_0 (
		.in({router_wrap_slice_IACK_2_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_0_ff_IACK_2_Q}),
		.sram(mux_tree_tapbuf_size2_409_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_409_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_409_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_2_1 (
		.in({router_wrap_slice_IACK_2_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_2_1_ff_IACK_2_Q}),
		.sram(mux_tree_tapbuf_size2_410_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_410_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_410_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_3_0 (
		.in({router_wrap_slice_IACK_3_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_0_ff_IACK_3_Q}),
		.sram(mux_tree_tapbuf_size2_411_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_411_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_411_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_3_1 (
		.in({router_wrap_slice_IACK_3_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_3_1_ff_IACK_3_Q}),
		.sram(mux_tree_tapbuf_size2_412_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_412_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_412_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_4_0 (
		.in({router_wrap_slice_IACK_4_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_0_ff_IACK_4_Q}),
		.sram(mux_tree_tapbuf_size2_413_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_413_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_413_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_IACK_4_1 (
		.in({router_wrap_slice_IACK_4_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_IACK_4_1_ff_IACK_4_Q}),
		.sram(mux_tree_tapbuf_size2_414_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_414_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_414_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_0_0 (
		.in({router_wrap_slice_ILCK_0_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_0_ff_ILCK_0_Q}),
		.sram(mux_tree_tapbuf_size2_415_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_415_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_415_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_0_1 (
		.in({router_wrap_slice_ILCK_0_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_0_1_ff_ILCK_0_Q}),
		.sram(mux_tree_tapbuf_size2_416_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_416_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_416_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_1_0 (
		.in({router_wrap_slice_ILCK_1_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_0_ff_ILCK_1_Q}),
		.sram(mux_tree_tapbuf_size2_417_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_417_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_417_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_1_1 (
		.in({router_wrap_slice_ILCK_1_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_1_1_ff_ILCK_1_Q}),
		.sram(mux_tree_tapbuf_size2_418_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_418_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_418_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_2_0 (
		.in({router_wrap_slice_ILCK_2_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_0_ff_ILCK_2_Q}),
		.sram(mux_tree_tapbuf_size2_419_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_419_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_419_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_2_1 (
		.in({router_wrap_slice_ILCK_2_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_2_1_ff_ILCK_2_Q}),
		.sram(mux_tree_tapbuf_size2_420_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_420_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_420_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_3_0 (
		.in({router_wrap_slice_ILCK_3_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_0_ff_ILCK_3_Q}),
		.sram(mux_tree_tapbuf_size2_421_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_421_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_421_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_3_1 (
		.in({router_wrap_slice_ILCK_3_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_3_1_ff_ILCK_3_Q}),
		.sram(mux_tree_tapbuf_size2_422_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_422_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_422_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_4_0 (
		.in({router_wrap_slice_ILCK_4_cfg[0], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_0_ff_ILCK_4_Q}),
		.sram(mux_tree_tapbuf_size2_423_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_423_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_423_out));

	mux_tree_tapbuf_size2 mux_router_wrap_0_ILCK_4_1 (
		.in({router_wrap_slice_ILCK_4_cfg[1], logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__ff_ILCK_4_1_ff_ILCK_4_Q}),
		.sram(mux_tree_tapbuf_size2_424_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_424_sram_inv[0:1]),
		.out(mux_tree_tapbuf_size2_424_out));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_0_cfg_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_1_cfg_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_82_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_83_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_84_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_85_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_86_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_87_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_88_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_89_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_90_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_91_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_92_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_93_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_94_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_95_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_96_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_97_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_98_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_99_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_100_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_101_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_102_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_103_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_2_cfg_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_104_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_105_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_106_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_107_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_108_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_109_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_110_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_111_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_112_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_113_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_114_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_115_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_116_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_117_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_118_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_119_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_120_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_121_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_122_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_123_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_124_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_125_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_126_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_127_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_128_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_129_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_130_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_131_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_132_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_133_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_134_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_135_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_136_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_137_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_137_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_138_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_138_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_3_cfg_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_139_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_139_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_140_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_140_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_141_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_141_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_142_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_142_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_143_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_143_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_144_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_144_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_145_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_145_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_146_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_146_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_147_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_147_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_148_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_148_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_149_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_149_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_150_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_150_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_151_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_151_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_152_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_152_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_153_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_153_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_154_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_154_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_155_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_155_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_156_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_156_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_157_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_157_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_158_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_158_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_159_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_159_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_160_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_160_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_161_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_161_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_162_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_162_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_163_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_163_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_164_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_164_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_165_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_165_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_166_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_166_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_167_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_167_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_168_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_168_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_169_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_169_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_170_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_170_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_171_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_171_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_172_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_172_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_173_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_173_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ODATA_4_cfg_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_174_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_174_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVALID_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_175_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_175_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVALID_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_176_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_176_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVALID_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_177_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_177_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVALID_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_178_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_178_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVALID_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_179_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_179_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVCH_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_180_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_180_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVCH_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_181_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_181_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVCH_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_182_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_182_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVCH_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_183_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_183_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OVCH_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_184_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_184_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_185_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_185_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_0_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_186_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_186_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_187_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_187_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_1_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_188_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_188_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_189_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_189_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_2_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_190_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_190_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_191_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_191_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_3_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_192_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_192_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_193_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_193_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OACK_4_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_194_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_194_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_195_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_195_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_0_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_196_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_196_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_197_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_197_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_1_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_198_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_198_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_199_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_199_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_2_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_200_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_200_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_201_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_201_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_3_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_202_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_202_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_203_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_203_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_ORDY_4_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_204_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_204_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_0_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_205_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_205_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_0_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_206_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_206_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_1_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_207_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_207_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_1_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_208_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_208_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_2_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_209_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_209_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_2_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_210_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_210_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_3_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_211_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_211_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_3_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_212_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_212_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_4_cfg_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_213_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_213_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_slice_OLCK_4_cfg_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_214_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_214_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_RST__0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_215_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_215_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_MY_XPOS_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_216_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_216_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_MY_XPOS_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_217_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_217_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_MY_YPOS_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_218_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_218_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_MY_YPOS_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_219_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_219_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_220_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_220_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_221_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_221_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_222_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_222_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_223_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_223_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_224_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_224_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_224_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_225_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_225_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_225_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_225_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_226_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_226_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_226_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_226_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_227_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_227_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_227_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_227_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_228_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_228_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_228_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_228_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_229_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_229_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_229_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_229_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_230_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_230_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_230_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_230_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_231_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_231_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_231_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_231_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_232_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_232_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_232_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_232_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_233_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_233_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_233_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_233_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_234_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_234_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_234_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_234_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_235_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_235_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_235_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_235_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_236_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_236_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_236_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_236_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_237_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_237_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_237_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_237_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_238_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_238_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_238_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_238_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_239_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_239_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_239_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_239_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_240_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_240_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_240_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_240_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_241_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_241_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_241_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_241_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_242_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_242_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_242_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_242_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_243_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_243_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_243_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_243_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_244_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_244_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_244_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_244_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_245_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_245_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_245_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_245_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_246_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_246_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_246_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_246_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_247_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_247_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_247_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_247_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_248_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_248_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_248_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_248_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_249_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_249_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_249_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_249_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_250_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_250_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_250_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_250_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_251_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_251_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_251_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_251_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_252_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_252_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_252_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_252_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_253_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_253_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_253_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_0_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_253_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_254_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_254_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_254_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_254_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_255_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_255_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_255_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_255_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_256_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_256_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_256_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_256_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_257_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_257_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_257_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_257_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_258_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_258_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_258_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_258_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_259_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_259_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_259_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_259_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_260_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_260_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_260_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_260_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_261_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_261_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_261_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_261_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_262_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_262_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_262_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_262_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_263_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_263_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_263_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_263_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_264_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_264_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_264_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_264_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_265_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_265_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_265_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_265_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_266_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_266_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_266_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_266_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_267_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_267_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_267_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_267_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_268_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_268_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_268_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_268_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_269_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_269_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_269_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_269_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_270_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_270_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_270_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_270_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_271_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_271_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_271_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_271_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_272_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_272_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_272_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_272_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_273_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_273_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_273_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_273_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_274_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_274_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_274_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_274_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_275_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_275_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_275_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_275_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_276_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_276_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_276_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_276_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_277_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_277_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_277_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_277_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_278_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_278_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_278_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_278_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_279_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_279_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_279_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_279_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_280_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_280_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_280_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_280_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_281_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_281_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_281_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_281_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_282_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_282_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_282_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_282_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_283_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_283_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_283_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_283_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_284_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_284_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_284_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_284_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_285_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_285_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_285_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_285_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_286_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_286_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_286_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_286_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_287_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_287_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_287_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_287_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_288_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_288_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_288_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_1_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_288_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_289_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_289_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_289_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_289_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_290_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_290_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_290_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_290_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_291_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_291_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_291_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_291_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_292_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_292_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_292_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_292_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_293_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_293_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_293_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_293_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_294_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_294_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_294_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_294_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_295_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_295_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_295_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_295_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_296_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_296_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_296_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_296_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_297_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_297_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_297_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_297_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_298_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_298_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_298_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_298_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_299_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_299_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_299_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_299_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_300_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_300_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_300_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_300_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_301_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_301_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_301_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_301_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_302_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_302_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_302_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_302_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_303_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_303_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_303_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_303_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_304_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_304_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_304_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_304_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_305_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_305_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_305_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_305_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_306_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_306_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_306_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_306_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_307_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_307_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_307_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_307_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_308_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_308_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_308_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_308_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_309_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_309_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_309_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_309_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_310_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_310_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_310_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_310_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_311_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_311_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_311_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_311_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_312_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_312_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_312_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_312_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_313_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_313_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_313_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_313_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_314_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_314_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_314_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_314_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_315_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_315_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_315_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_315_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_316_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_316_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_316_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_316_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_317_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_317_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_317_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_317_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_318_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_318_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_318_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_318_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_319_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_319_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_319_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_319_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_320_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_320_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_320_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_320_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_321_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_321_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_321_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_321_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_322_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_322_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_322_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_322_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_323_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_323_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_323_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_2_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_323_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_324_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_324_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_324_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_324_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_325_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_325_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_325_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_325_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_326_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_326_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_326_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_326_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_327_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_327_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_327_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_327_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_328_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_328_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_328_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_328_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_329_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_329_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_329_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_329_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_330_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_330_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_330_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_330_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_331_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_331_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_331_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_331_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_332_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_332_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_332_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_332_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_333_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_333_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_333_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_333_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_334_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_334_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_334_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_334_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_335_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_335_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_335_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_335_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_336_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_336_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_336_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_336_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_337_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_337_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_337_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_337_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_338_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_338_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_338_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_338_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_339_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_339_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_339_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_339_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_340_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_340_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_340_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_340_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_341_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_341_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_341_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_341_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_342_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_342_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_342_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_342_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_343_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_343_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_343_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_343_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_344_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_344_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_344_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_344_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_345_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_345_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_345_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_345_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_346_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_346_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_346_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_346_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_347_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_347_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_347_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_347_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_348_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_348_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_348_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_348_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_349_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_349_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_349_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_349_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_350_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_350_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_350_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_350_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_351_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_351_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_351_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_351_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_352_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_352_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_352_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_352_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_353_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_353_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_353_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_353_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_354_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_354_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_354_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_354_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_355_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_355_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_355_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_355_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_356_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_356_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_356_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_356_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_357_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_357_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_357_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_357_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_358_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_358_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_358_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_3_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_358_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_359_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_359_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_359_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_359_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_360_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_360_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_360_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_360_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_361_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_361_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_361_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_361_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_362_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_362_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_362_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_362_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_363_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_363_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_363_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_363_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_364_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_364_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_364_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_364_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_365_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_365_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_365_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_365_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_366_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_366_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_366_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_366_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_367_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_367_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_367_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_367_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_368_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_368_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_368_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_368_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_369_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_369_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_369_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_369_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_370_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_370_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_370_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_370_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_371_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_371_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_371_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_371_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_372_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_372_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_372_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_372_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_373_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_373_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_373_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_373_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_374_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_374_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_374_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_374_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_375_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_375_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_375_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_375_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_376_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_376_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_376_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_376_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_377_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_377_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_377_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_377_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_378_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_378_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_378_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_378_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_379_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_379_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_379_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_379_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_380_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_380_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_380_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_380_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_381_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_381_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_381_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_381_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_382_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_382_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_382_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_382_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_383_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_383_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_383_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_383_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_384_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_384_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_384_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_384_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_385_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_385_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_385_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_385_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_386_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_386_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_386_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_386_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_387_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_387_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_387_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_387_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_388_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_388_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_388_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_388_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_389_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_389_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_389_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_389_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_390_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_390_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_390_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_390_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_391_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_391_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_391_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_391_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_392_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_392_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_392_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_392_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_393_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_393_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_393_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IDATA_4_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_393_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_394_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_394_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_394_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVALID_0_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_394_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_395_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_395_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_395_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVALID_1_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_395_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_396_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_396_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_396_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVALID_2_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_396_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_397_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_397_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_397_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVALID_3_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_397_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_398_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_398_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_398_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVALID_4_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_398_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_399_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_399_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_399_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVCH_0_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_399_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_400_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_400_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_400_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVCH_1_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_400_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_401_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_401_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_401_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVCH_2_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_401_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_402_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_402_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_402_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVCH_3_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_402_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_403_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_403_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_403_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IVCH_4_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_403_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_404_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_404_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_404_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_0_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_404_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_405_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_405_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_405_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_0_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_405_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_406_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_406_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_406_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_1_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_406_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_407_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_407_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_407_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_1_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_407_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_408_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_408_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_408_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_2_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_408_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_409_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_409_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_409_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_2_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_409_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_410_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_410_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_410_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_3_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_410_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_411_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_411_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_411_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_3_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_411_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_412_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_412_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_412_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_4_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_412_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_413_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_413_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_413_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_IACK_4_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_413_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_414_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_414_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_414_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_0_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_414_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_415_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_415_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_415_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_0_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_415_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_416_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_416_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_416_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_1_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_416_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_417_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_417_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_417_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_1_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_417_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_418_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_418_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_418_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_2_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_418_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_419_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_419_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_419_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_2_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_419_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_420_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_420_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_420_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_3_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_420_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_421_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_421_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_421_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_3_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_421_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_422_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_422_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_422_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_4_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_422_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_423_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_423_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_423_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_router_wrap_0_ILCK_4_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_423_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_424_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_424_sram_inv[0:1]));

	direct_interc direct_interc_0_ (
		.in(router_wrap_slice_RST__cfg),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(router_wrap_slice_MY_XPOS_cfg[0]),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(router_wrap_slice_MY_XPOS_cfg[1]),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(router_wrap_slice_MY_YPOS_cfg[0]),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(router_wrap_slice_MY_YPOS_cfg[1]),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(router_wrap_slice_IDATA_0_cfg[0]),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(router_wrap_slice_IDATA_0_cfg[1]),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(router_wrap_slice_IDATA_0_cfg[2]),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(router_wrap_slice_IDATA_0_cfg[3]),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(router_wrap_slice_IDATA_0_cfg[4]),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(router_wrap_slice_IDATA_0_cfg[5]),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(router_wrap_slice_IDATA_0_cfg[6]),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(router_wrap_slice_IDATA_0_cfg[7]),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(router_wrap_slice_IDATA_0_cfg[8]),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(router_wrap_slice_IDATA_0_cfg[9]),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_29_out));

	direct_interc direct_interc_30_ (
		.in(router_wrap_slice_IDATA_0_cfg[10]),
		.out(direct_interc_30_out));

	direct_interc direct_interc_31_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_31_out));

	direct_interc direct_interc_32_ (
		.in(router_wrap_slice_IDATA_0_cfg[11]),
		.out(direct_interc_32_out));

	direct_interc direct_interc_33_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_33_out));

	direct_interc direct_interc_34_ (
		.in(router_wrap_slice_IDATA_0_cfg[12]),
		.out(direct_interc_34_out));

	direct_interc direct_interc_35_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_35_out));

	direct_interc direct_interc_36_ (
		.in(router_wrap_slice_IDATA_0_cfg[13]),
		.out(direct_interc_36_out));

	direct_interc direct_interc_37_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_37_out));

	direct_interc direct_interc_38_ (
		.in(router_wrap_slice_IDATA_0_cfg[14]),
		.out(direct_interc_38_out));

	direct_interc direct_interc_39_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_39_out));

	direct_interc direct_interc_40_ (
		.in(router_wrap_slice_IDATA_0_cfg[15]),
		.out(direct_interc_40_out));

	direct_interc direct_interc_41_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_41_out));

	direct_interc direct_interc_42_ (
		.in(router_wrap_slice_IDATA_0_cfg[16]),
		.out(direct_interc_42_out));

	direct_interc direct_interc_43_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_43_out));

	direct_interc direct_interc_44_ (
		.in(router_wrap_slice_IDATA_0_cfg[17]),
		.out(direct_interc_44_out));

	direct_interc direct_interc_45_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_45_out));

	direct_interc direct_interc_46_ (
		.in(router_wrap_slice_IDATA_0_cfg[18]),
		.out(direct_interc_46_out));

	direct_interc direct_interc_47_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_47_out));

	direct_interc direct_interc_48_ (
		.in(router_wrap_slice_IDATA_0_cfg[19]),
		.out(direct_interc_48_out));

	direct_interc direct_interc_49_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_49_out));

	direct_interc direct_interc_50_ (
		.in(router_wrap_slice_IDATA_0_cfg[20]),
		.out(direct_interc_50_out));

	direct_interc direct_interc_51_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_51_out));

	direct_interc direct_interc_52_ (
		.in(router_wrap_slice_IDATA_0_cfg[21]),
		.out(direct_interc_52_out));

	direct_interc direct_interc_53_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_53_out));

	direct_interc direct_interc_54_ (
		.in(router_wrap_slice_IDATA_0_cfg[22]),
		.out(direct_interc_54_out));

	direct_interc direct_interc_55_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_55_out));

	direct_interc direct_interc_56_ (
		.in(router_wrap_slice_IDATA_0_cfg[23]),
		.out(direct_interc_56_out));

	direct_interc direct_interc_57_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_57_out));

	direct_interc direct_interc_58_ (
		.in(router_wrap_slice_IDATA_0_cfg[24]),
		.out(direct_interc_58_out));

	direct_interc direct_interc_59_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_59_out));

	direct_interc direct_interc_60_ (
		.in(router_wrap_slice_IDATA_0_cfg[25]),
		.out(direct_interc_60_out));

	direct_interc direct_interc_61_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_61_out));

	direct_interc direct_interc_62_ (
		.in(router_wrap_slice_IDATA_0_cfg[26]),
		.out(direct_interc_62_out));

	direct_interc direct_interc_63_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_63_out));

	direct_interc direct_interc_64_ (
		.in(router_wrap_slice_IDATA_0_cfg[27]),
		.out(direct_interc_64_out));

	direct_interc direct_interc_65_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_65_out));

	direct_interc direct_interc_66_ (
		.in(router_wrap_slice_IDATA_0_cfg[28]),
		.out(direct_interc_66_out));

	direct_interc direct_interc_67_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_67_out));

	direct_interc direct_interc_68_ (
		.in(router_wrap_slice_IDATA_0_cfg[29]),
		.out(direct_interc_68_out));

	direct_interc direct_interc_69_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_69_out));

	direct_interc direct_interc_70_ (
		.in(router_wrap_slice_IDATA_0_cfg[30]),
		.out(direct_interc_70_out));

	direct_interc direct_interc_71_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_71_out));

	direct_interc direct_interc_72_ (
		.in(router_wrap_slice_IDATA_0_cfg[31]),
		.out(direct_interc_72_out));

	direct_interc direct_interc_73_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_73_out));

	direct_interc direct_interc_74_ (
		.in(router_wrap_slice_IDATA_0_cfg[32]),
		.out(direct_interc_74_out));

	direct_interc direct_interc_75_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_75_out));

	direct_interc direct_interc_76_ (
		.in(router_wrap_slice_IDATA_0_cfg[33]),
		.out(direct_interc_76_out));

	direct_interc direct_interc_77_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_77_out));

	direct_interc direct_interc_78_ (
		.in(router_wrap_slice_IDATA_0_cfg[34]),
		.out(direct_interc_78_out));

	direct_interc direct_interc_79_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_79_out));

	direct_interc direct_interc_80_ (
		.in(router_wrap_slice_IDATA_1_cfg[0]),
		.out(direct_interc_80_out));

	direct_interc direct_interc_81_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_81_out));

	direct_interc direct_interc_82_ (
		.in(router_wrap_slice_IDATA_1_cfg[1]),
		.out(direct_interc_82_out));

	direct_interc direct_interc_83_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_83_out));

	direct_interc direct_interc_84_ (
		.in(router_wrap_slice_IDATA_1_cfg[2]),
		.out(direct_interc_84_out));

	direct_interc direct_interc_85_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_85_out));

	direct_interc direct_interc_86_ (
		.in(router_wrap_slice_IDATA_1_cfg[3]),
		.out(direct_interc_86_out));

	direct_interc direct_interc_87_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_87_out));

	direct_interc direct_interc_88_ (
		.in(router_wrap_slice_IDATA_1_cfg[4]),
		.out(direct_interc_88_out));

	direct_interc direct_interc_89_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_89_out));

	direct_interc direct_interc_90_ (
		.in(router_wrap_slice_IDATA_1_cfg[5]),
		.out(direct_interc_90_out));

	direct_interc direct_interc_91_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_91_out));

	direct_interc direct_interc_92_ (
		.in(router_wrap_slice_IDATA_1_cfg[6]),
		.out(direct_interc_92_out));

	direct_interc direct_interc_93_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_93_out));

	direct_interc direct_interc_94_ (
		.in(router_wrap_slice_IDATA_1_cfg[7]),
		.out(direct_interc_94_out));

	direct_interc direct_interc_95_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_95_out));

	direct_interc direct_interc_96_ (
		.in(router_wrap_slice_IDATA_1_cfg[8]),
		.out(direct_interc_96_out));

	direct_interc direct_interc_97_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_97_out));

	direct_interc direct_interc_98_ (
		.in(router_wrap_slice_IDATA_1_cfg[9]),
		.out(direct_interc_98_out));

	direct_interc direct_interc_99_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_99_out));

	direct_interc direct_interc_100_ (
		.in(router_wrap_slice_IDATA_1_cfg[10]),
		.out(direct_interc_100_out));

	direct_interc direct_interc_101_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_101_out));

	direct_interc direct_interc_102_ (
		.in(router_wrap_slice_IDATA_1_cfg[11]),
		.out(direct_interc_102_out));

	direct_interc direct_interc_103_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_103_out));

	direct_interc direct_interc_104_ (
		.in(router_wrap_slice_IDATA_1_cfg[12]),
		.out(direct_interc_104_out));

	direct_interc direct_interc_105_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_105_out));

	direct_interc direct_interc_106_ (
		.in(router_wrap_slice_IDATA_1_cfg[13]),
		.out(direct_interc_106_out));

	direct_interc direct_interc_107_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_107_out));

	direct_interc direct_interc_108_ (
		.in(router_wrap_slice_IDATA_1_cfg[14]),
		.out(direct_interc_108_out));

	direct_interc direct_interc_109_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_109_out));

	direct_interc direct_interc_110_ (
		.in(router_wrap_slice_IDATA_1_cfg[15]),
		.out(direct_interc_110_out));

	direct_interc direct_interc_111_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_111_out));

	direct_interc direct_interc_112_ (
		.in(router_wrap_slice_IDATA_1_cfg[16]),
		.out(direct_interc_112_out));

	direct_interc direct_interc_113_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_113_out));

	direct_interc direct_interc_114_ (
		.in(router_wrap_slice_IDATA_1_cfg[17]),
		.out(direct_interc_114_out));

	direct_interc direct_interc_115_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_115_out));

	direct_interc direct_interc_116_ (
		.in(router_wrap_slice_IDATA_1_cfg[18]),
		.out(direct_interc_116_out));

	direct_interc direct_interc_117_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_117_out));

	direct_interc direct_interc_118_ (
		.in(router_wrap_slice_IDATA_1_cfg[19]),
		.out(direct_interc_118_out));

	direct_interc direct_interc_119_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_119_out));

	direct_interc direct_interc_120_ (
		.in(router_wrap_slice_IDATA_1_cfg[20]),
		.out(direct_interc_120_out));

	direct_interc direct_interc_121_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_121_out));

	direct_interc direct_interc_122_ (
		.in(router_wrap_slice_IDATA_1_cfg[21]),
		.out(direct_interc_122_out));

	direct_interc direct_interc_123_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_123_out));

	direct_interc direct_interc_124_ (
		.in(router_wrap_slice_IDATA_1_cfg[22]),
		.out(direct_interc_124_out));

	direct_interc direct_interc_125_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_125_out));

	direct_interc direct_interc_126_ (
		.in(router_wrap_slice_IDATA_1_cfg[23]),
		.out(direct_interc_126_out));

	direct_interc direct_interc_127_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_127_out));

	direct_interc direct_interc_128_ (
		.in(router_wrap_slice_IDATA_1_cfg[24]),
		.out(direct_interc_128_out));

	direct_interc direct_interc_129_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_129_out));

	direct_interc direct_interc_130_ (
		.in(router_wrap_slice_IDATA_1_cfg[25]),
		.out(direct_interc_130_out));

	direct_interc direct_interc_131_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_131_out));

	direct_interc direct_interc_132_ (
		.in(router_wrap_slice_IDATA_1_cfg[26]),
		.out(direct_interc_132_out));

	direct_interc direct_interc_133_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_133_out));

	direct_interc direct_interc_134_ (
		.in(router_wrap_slice_IDATA_1_cfg[27]),
		.out(direct_interc_134_out));

	direct_interc direct_interc_135_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_135_out));

	direct_interc direct_interc_136_ (
		.in(router_wrap_slice_IDATA_1_cfg[28]),
		.out(direct_interc_136_out));

	direct_interc direct_interc_137_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_137_out));

	direct_interc direct_interc_138_ (
		.in(router_wrap_slice_IDATA_1_cfg[29]),
		.out(direct_interc_138_out));

	direct_interc direct_interc_139_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_139_out));

	direct_interc direct_interc_140_ (
		.in(router_wrap_slice_IDATA_1_cfg[30]),
		.out(direct_interc_140_out));

	direct_interc direct_interc_141_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_141_out));

	direct_interc direct_interc_142_ (
		.in(router_wrap_slice_IDATA_1_cfg[31]),
		.out(direct_interc_142_out));

	direct_interc direct_interc_143_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_143_out));

	direct_interc direct_interc_144_ (
		.in(router_wrap_slice_IDATA_1_cfg[32]),
		.out(direct_interc_144_out));

	direct_interc direct_interc_145_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_145_out));

	direct_interc direct_interc_146_ (
		.in(router_wrap_slice_IDATA_1_cfg[33]),
		.out(direct_interc_146_out));

	direct_interc direct_interc_147_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_147_out));

	direct_interc direct_interc_148_ (
		.in(router_wrap_slice_IDATA_1_cfg[34]),
		.out(direct_interc_148_out));

	direct_interc direct_interc_149_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_149_out));

	direct_interc direct_interc_150_ (
		.in(router_wrap_slice_IDATA_2_cfg[0]),
		.out(direct_interc_150_out));

	direct_interc direct_interc_151_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_151_out));

	direct_interc direct_interc_152_ (
		.in(router_wrap_slice_IDATA_2_cfg[1]),
		.out(direct_interc_152_out));

	direct_interc direct_interc_153_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_153_out));

	direct_interc direct_interc_154_ (
		.in(router_wrap_slice_IDATA_2_cfg[2]),
		.out(direct_interc_154_out));

	direct_interc direct_interc_155_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_155_out));

	direct_interc direct_interc_156_ (
		.in(router_wrap_slice_IDATA_2_cfg[3]),
		.out(direct_interc_156_out));

	direct_interc direct_interc_157_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_157_out));

	direct_interc direct_interc_158_ (
		.in(router_wrap_slice_IDATA_2_cfg[4]),
		.out(direct_interc_158_out));

	direct_interc direct_interc_159_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_159_out));

	direct_interc direct_interc_160_ (
		.in(router_wrap_slice_IDATA_2_cfg[5]),
		.out(direct_interc_160_out));

	direct_interc direct_interc_161_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_161_out));

	direct_interc direct_interc_162_ (
		.in(router_wrap_slice_IDATA_2_cfg[6]),
		.out(direct_interc_162_out));

	direct_interc direct_interc_163_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_163_out));

	direct_interc direct_interc_164_ (
		.in(router_wrap_slice_IDATA_2_cfg[7]),
		.out(direct_interc_164_out));

	direct_interc direct_interc_165_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_165_out));

	direct_interc direct_interc_166_ (
		.in(router_wrap_slice_IDATA_2_cfg[8]),
		.out(direct_interc_166_out));

	direct_interc direct_interc_167_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_167_out));

	direct_interc direct_interc_168_ (
		.in(router_wrap_slice_IDATA_2_cfg[9]),
		.out(direct_interc_168_out));

	direct_interc direct_interc_169_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_169_out));

	direct_interc direct_interc_170_ (
		.in(router_wrap_slice_IDATA_2_cfg[10]),
		.out(direct_interc_170_out));

	direct_interc direct_interc_171_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_171_out));

	direct_interc direct_interc_172_ (
		.in(router_wrap_slice_IDATA_2_cfg[11]),
		.out(direct_interc_172_out));

	direct_interc direct_interc_173_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_173_out));

	direct_interc direct_interc_174_ (
		.in(router_wrap_slice_IDATA_2_cfg[12]),
		.out(direct_interc_174_out));

	direct_interc direct_interc_175_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_175_out));

	direct_interc direct_interc_176_ (
		.in(router_wrap_slice_IDATA_2_cfg[13]),
		.out(direct_interc_176_out));

	direct_interc direct_interc_177_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_177_out));

	direct_interc direct_interc_178_ (
		.in(router_wrap_slice_IDATA_2_cfg[14]),
		.out(direct_interc_178_out));

	direct_interc direct_interc_179_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_179_out));

	direct_interc direct_interc_180_ (
		.in(router_wrap_slice_IDATA_2_cfg[15]),
		.out(direct_interc_180_out));

	direct_interc direct_interc_181_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_181_out));

	direct_interc direct_interc_182_ (
		.in(router_wrap_slice_IDATA_2_cfg[16]),
		.out(direct_interc_182_out));

	direct_interc direct_interc_183_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_183_out));

	direct_interc direct_interc_184_ (
		.in(router_wrap_slice_IDATA_2_cfg[17]),
		.out(direct_interc_184_out));

	direct_interc direct_interc_185_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_185_out));

	direct_interc direct_interc_186_ (
		.in(router_wrap_slice_IDATA_2_cfg[18]),
		.out(direct_interc_186_out));

	direct_interc direct_interc_187_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_187_out));

	direct_interc direct_interc_188_ (
		.in(router_wrap_slice_IDATA_2_cfg[19]),
		.out(direct_interc_188_out));

	direct_interc direct_interc_189_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_189_out));

	direct_interc direct_interc_190_ (
		.in(router_wrap_slice_IDATA_2_cfg[20]),
		.out(direct_interc_190_out));

	direct_interc direct_interc_191_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_191_out));

	direct_interc direct_interc_192_ (
		.in(router_wrap_slice_IDATA_2_cfg[21]),
		.out(direct_interc_192_out));

	direct_interc direct_interc_193_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_193_out));

	direct_interc direct_interc_194_ (
		.in(router_wrap_slice_IDATA_2_cfg[22]),
		.out(direct_interc_194_out));

	direct_interc direct_interc_195_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_195_out));

	direct_interc direct_interc_196_ (
		.in(router_wrap_slice_IDATA_2_cfg[23]),
		.out(direct_interc_196_out));

	direct_interc direct_interc_197_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_197_out));

	direct_interc direct_interc_198_ (
		.in(router_wrap_slice_IDATA_2_cfg[24]),
		.out(direct_interc_198_out));

	direct_interc direct_interc_199_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_199_out));

	direct_interc direct_interc_200_ (
		.in(router_wrap_slice_IDATA_2_cfg[25]),
		.out(direct_interc_200_out));

	direct_interc direct_interc_201_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_201_out));

	direct_interc direct_interc_202_ (
		.in(router_wrap_slice_IDATA_2_cfg[26]),
		.out(direct_interc_202_out));

	direct_interc direct_interc_203_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_203_out));

	direct_interc direct_interc_204_ (
		.in(router_wrap_slice_IDATA_2_cfg[27]),
		.out(direct_interc_204_out));

	direct_interc direct_interc_205_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_205_out));

	direct_interc direct_interc_206_ (
		.in(router_wrap_slice_IDATA_2_cfg[28]),
		.out(direct_interc_206_out));

	direct_interc direct_interc_207_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_207_out));

	direct_interc direct_interc_208_ (
		.in(router_wrap_slice_IDATA_2_cfg[29]),
		.out(direct_interc_208_out));

	direct_interc direct_interc_209_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_209_out));

	direct_interc direct_interc_210_ (
		.in(router_wrap_slice_IDATA_2_cfg[30]),
		.out(direct_interc_210_out));

	direct_interc direct_interc_211_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_211_out));

	direct_interc direct_interc_212_ (
		.in(router_wrap_slice_IDATA_2_cfg[31]),
		.out(direct_interc_212_out));

	direct_interc direct_interc_213_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_213_out));

	direct_interc direct_interc_214_ (
		.in(router_wrap_slice_IDATA_2_cfg[32]),
		.out(direct_interc_214_out));

	direct_interc direct_interc_215_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_215_out));

	direct_interc direct_interc_216_ (
		.in(router_wrap_slice_IDATA_2_cfg[33]),
		.out(direct_interc_216_out));

	direct_interc direct_interc_217_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_217_out));

	direct_interc direct_interc_218_ (
		.in(router_wrap_slice_IDATA_2_cfg[34]),
		.out(direct_interc_218_out));

	direct_interc direct_interc_219_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_219_out));

	direct_interc direct_interc_220_ (
		.in(router_wrap_slice_IDATA_3_cfg[0]),
		.out(direct_interc_220_out));

	direct_interc direct_interc_221_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_221_out));

	direct_interc direct_interc_222_ (
		.in(router_wrap_slice_IDATA_3_cfg[1]),
		.out(direct_interc_222_out));

	direct_interc direct_interc_223_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_223_out));

	direct_interc direct_interc_224_ (
		.in(router_wrap_slice_IDATA_3_cfg[2]),
		.out(direct_interc_224_out));

	direct_interc direct_interc_225_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_225_out));

	direct_interc direct_interc_226_ (
		.in(router_wrap_slice_IDATA_3_cfg[3]),
		.out(direct_interc_226_out));

	direct_interc direct_interc_227_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_227_out));

	direct_interc direct_interc_228_ (
		.in(router_wrap_slice_IDATA_3_cfg[4]),
		.out(direct_interc_228_out));

	direct_interc direct_interc_229_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_229_out));

	direct_interc direct_interc_230_ (
		.in(router_wrap_slice_IDATA_3_cfg[5]),
		.out(direct_interc_230_out));

	direct_interc direct_interc_231_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_231_out));

	direct_interc direct_interc_232_ (
		.in(router_wrap_slice_IDATA_3_cfg[6]),
		.out(direct_interc_232_out));

	direct_interc direct_interc_233_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_233_out));

	direct_interc direct_interc_234_ (
		.in(router_wrap_slice_IDATA_3_cfg[7]),
		.out(direct_interc_234_out));

	direct_interc direct_interc_235_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_235_out));

	direct_interc direct_interc_236_ (
		.in(router_wrap_slice_IDATA_3_cfg[8]),
		.out(direct_interc_236_out));

	direct_interc direct_interc_237_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_237_out));

	direct_interc direct_interc_238_ (
		.in(router_wrap_slice_IDATA_3_cfg[9]),
		.out(direct_interc_238_out));

	direct_interc direct_interc_239_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_239_out));

	direct_interc direct_interc_240_ (
		.in(router_wrap_slice_IDATA_3_cfg[10]),
		.out(direct_interc_240_out));

	direct_interc direct_interc_241_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_241_out));

	direct_interc direct_interc_242_ (
		.in(router_wrap_slice_IDATA_3_cfg[11]),
		.out(direct_interc_242_out));

	direct_interc direct_interc_243_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_243_out));

	direct_interc direct_interc_244_ (
		.in(router_wrap_slice_IDATA_3_cfg[12]),
		.out(direct_interc_244_out));

	direct_interc direct_interc_245_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_245_out));

	direct_interc direct_interc_246_ (
		.in(router_wrap_slice_IDATA_3_cfg[13]),
		.out(direct_interc_246_out));

	direct_interc direct_interc_247_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_247_out));

	direct_interc direct_interc_248_ (
		.in(router_wrap_slice_IDATA_3_cfg[14]),
		.out(direct_interc_248_out));

	direct_interc direct_interc_249_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_249_out));

	direct_interc direct_interc_250_ (
		.in(router_wrap_slice_IDATA_3_cfg[15]),
		.out(direct_interc_250_out));

	direct_interc direct_interc_251_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_251_out));

	direct_interc direct_interc_252_ (
		.in(router_wrap_slice_IDATA_3_cfg[16]),
		.out(direct_interc_252_out));

	direct_interc direct_interc_253_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_253_out));

	direct_interc direct_interc_254_ (
		.in(router_wrap_slice_IDATA_3_cfg[17]),
		.out(direct_interc_254_out));

	direct_interc direct_interc_255_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_255_out));

	direct_interc direct_interc_256_ (
		.in(router_wrap_slice_IDATA_3_cfg[18]),
		.out(direct_interc_256_out));

	direct_interc direct_interc_257_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_257_out));

	direct_interc direct_interc_258_ (
		.in(router_wrap_slice_IDATA_3_cfg[19]),
		.out(direct_interc_258_out));

	direct_interc direct_interc_259_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_259_out));

	direct_interc direct_interc_260_ (
		.in(router_wrap_slice_IDATA_3_cfg[20]),
		.out(direct_interc_260_out));

	direct_interc direct_interc_261_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_261_out));

	direct_interc direct_interc_262_ (
		.in(router_wrap_slice_IDATA_3_cfg[21]),
		.out(direct_interc_262_out));

	direct_interc direct_interc_263_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_263_out));

	direct_interc direct_interc_264_ (
		.in(router_wrap_slice_IDATA_3_cfg[22]),
		.out(direct_interc_264_out));

	direct_interc direct_interc_265_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_265_out));

	direct_interc direct_interc_266_ (
		.in(router_wrap_slice_IDATA_3_cfg[23]),
		.out(direct_interc_266_out));

	direct_interc direct_interc_267_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_267_out));

	direct_interc direct_interc_268_ (
		.in(router_wrap_slice_IDATA_3_cfg[24]),
		.out(direct_interc_268_out));

	direct_interc direct_interc_269_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_269_out));

	direct_interc direct_interc_270_ (
		.in(router_wrap_slice_IDATA_3_cfg[25]),
		.out(direct_interc_270_out));

	direct_interc direct_interc_271_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_271_out));

	direct_interc direct_interc_272_ (
		.in(router_wrap_slice_IDATA_3_cfg[26]),
		.out(direct_interc_272_out));

	direct_interc direct_interc_273_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_273_out));

	direct_interc direct_interc_274_ (
		.in(router_wrap_slice_IDATA_3_cfg[27]),
		.out(direct_interc_274_out));

	direct_interc direct_interc_275_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_275_out));

	direct_interc direct_interc_276_ (
		.in(router_wrap_slice_IDATA_3_cfg[28]),
		.out(direct_interc_276_out));

	direct_interc direct_interc_277_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_277_out));

	direct_interc direct_interc_278_ (
		.in(router_wrap_slice_IDATA_3_cfg[29]),
		.out(direct_interc_278_out));

	direct_interc direct_interc_279_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_279_out));

	direct_interc direct_interc_280_ (
		.in(router_wrap_slice_IDATA_3_cfg[30]),
		.out(direct_interc_280_out));

	direct_interc direct_interc_281_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_281_out));

	direct_interc direct_interc_282_ (
		.in(router_wrap_slice_IDATA_3_cfg[31]),
		.out(direct_interc_282_out));

	direct_interc direct_interc_283_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_283_out));

	direct_interc direct_interc_284_ (
		.in(router_wrap_slice_IDATA_3_cfg[32]),
		.out(direct_interc_284_out));

	direct_interc direct_interc_285_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_285_out));

	direct_interc direct_interc_286_ (
		.in(router_wrap_slice_IDATA_3_cfg[33]),
		.out(direct_interc_286_out));

	direct_interc direct_interc_287_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_287_out));

	direct_interc direct_interc_288_ (
		.in(router_wrap_slice_IDATA_3_cfg[34]),
		.out(direct_interc_288_out));

	direct_interc direct_interc_289_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_289_out));

	direct_interc direct_interc_290_ (
		.in(router_wrap_slice_IDATA_4_cfg[0]),
		.out(direct_interc_290_out));

	direct_interc direct_interc_291_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_291_out));

	direct_interc direct_interc_292_ (
		.in(router_wrap_slice_IDATA_4_cfg[1]),
		.out(direct_interc_292_out));

	direct_interc direct_interc_293_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_293_out));

	direct_interc direct_interc_294_ (
		.in(router_wrap_slice_IDATA_4_cfg[2]),
		.out(direct_interc_294_out));

	direct_interc direct_interc_295_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_295_out));

	direct_interc direct_interc_296_ (
		.in(router_wrap_slice_IDATA_4_cfg[3]),
		.out(direct_interc_296_out));

	direct_interc direct_interc_297_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_297_out));

	direct_interc direct_interc_298_ (
		.in(router_wrap_slice_IDATA_4_cfg[4]),
		.out(direct_interc_298_out));

	direct_interc direct_interc_299_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_299_out));

	direct_interc direct_interc_300_ (
		.in(router_wrap_slice_IDATA_4_cfg[5]),
		.out(direct_interc_300_out));

	direct_interc direct_interc_301_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_301_out));

	direct_interc direct_interc_302_ (
		.in(router_wrap_slice_IDATA_4_cfg[6]),
		.out(direct_interc_302_out));

	direct_interc direct_interc_303_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_303_out));

	direct_interc direct_interc_304_ (
		.in(router_wrap_slice_IDATA_4_cfg[7]),
		.out(direct_interc_304_out));

	direct_interc direct_interc_305_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_305_out));

	direct_interc direct_interc_306_ (
		.in(router_wrap_slice_IDATA_4_cfg[8]),
		.out(direct_interc_306_out));

	direct_interc direct_interc_307_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_307_out));

	direct_interc direct_interc_308_ (
		.in(router_wrap_slice_IDATA_4_cfg[9]),
		.out(direct_interc_308_out));

	direct_interc direct_interc_309_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_309_out));

	direct_interc direct_interc_310_ (
		.in(router_wrap_slice_IDATA_4_cfg[10]),
		.out(direct_interc_310_out));

	direct_interc direct_interc_311_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_311_out));

	direct_interc direct_interc_312_ (
		.in(router_wrap_slice_IDATA_4_cfg[11]),
		.out(direct_interc_312_out));

	direct_interc direct_interc_313_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_313_out));

	direct_interc direct_interc_314_ (
		.in(router_wrap_slice_IDATA_4_cfg[12]),
		.out(direct_interc_314_out));

	direct_interc direct_interc_315_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_315_out));

	direct_interc direct_interc_316_ (
		.in(router_wrap_slice_IDATA_4_cfg[13]),
		.out(direct_interc_316_out));

	direct_interc direct_interc_317_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_317_out));

	direct_interc direct_interc_318_ (
		.in(router_wrap_slice_IDATA_4_cfg[14]),
		.out(direct_interc_318_out));

	direct_interc direct_interc_319_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_319_out));

	direct_interc direct_interc_320_ (
		.in(router_wrap_slice_IDATA_4_cfg[15]),
		.out(direct_interc_320_out));

	direct_interc direct_interc_321_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_321_out));

	direct_interc direct_interc_322_ (
		.in(router_wrap_slice_IDATA_4_cfg[16]),
		.out(direct_interc_322_out));

	direct_interc direct_interc_323_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_323_out));

	direct_interc direct_interc_324_ (
		.in(router_wrap_slice_IDATA_4_cfg[17]),
		.out(direct_interc_324_out));

	direct_interc direct_interc_325_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_325_out));

	direct_interc direct_interc_326_ (
		.in(router_wrap_slice_IDATA_4_cfg[18]),
		.out(direct_interc_326_out));

	direct_interc direct_interc_327_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_327_out));

	direct_interc direct_interc_328_ (
		.in(router_wrap_slice_IDATA_4_cfg[19]),
		.out(direct_interc_328_out));

	direct_interc direct_interc_329_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_329_out));

	direct_interc direct_interc_330_ (
		.in(router_wrap_slice_IDATA_4_cfg[20]),
		.out(direct_interc_330_out));

	direct_interc direct_interc_331_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_331_out));

	direct_interc direct_interc_332_ (
		.in(router_wrap_slice_IDATA_4_cfg[21]),
		.out(direct_interc_332_out));

	direct_interc direct_interc_333_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_333_out));

	direct_interc direct_interc_334_ (
		.in(router_wrap_slice_IDATA_4_cfg[22]),
		.out(direct_interc_334_out));

	direct_interc direct_interc_335_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_335_out));

	direct_interc direct_interc_336_ (
		.in(router_wrap_slice_IDATA_4_cfg[23]),
		.out(direct_interc_336_out));

	direct_interc direct_interc_337_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_337_out));

	direct_interc direct_interc_338_ (
		.in(router_wrap_slice_IDATA_4_cfg[24]),
		.out(direct_interc_338_out));

	direct_interc direct_interc_339_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_339_out));

	direct_interc direct_interc_340_ (
		.in(router_wrap_slice_IDATA_4_cfg[25]),
		.out(direct_interc_340_out));

	direct_interc direct_interc_341_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_341_out));

	direct_interc direct_interc_342_ (
		.in(router_wrap_slice_IDATA_4_cfg[26]),
		.out(direct_interc_342_out));

	direct_interc direct_interc_343_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_343_out));

	direct_interc direct_interc_344_ (
		.in(router_wrap_slice_IDATA_4_cfg[27]),
		.out(direct_interc_344_out));

	direct_interc direct_interc_345_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_345_out));

	direct_interc direct_interc_346_ (
		.in(router_wrap_slice_IDATA_4_cfg[28]),
		.out(direct_interc_346_out));

	direct_interc direct_interc_347_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_347_out));

	direct_interc direct_interc_348_ (
		.in(router_wrap_slice_IDATA_4_cfg[29]),
		.out(direct_interc_348_out));

	direct_interc direct_interc_349_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_349_out));

	direct_interc direct_interc_350_ (
		.in(router_wrap_slice_IDATA_4_cfg[30]),
		.out(direct_interc_350_out));

	direct_interc direct_interc_351_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_351_out));

	direct_interc direct_interc_352_ (
		.in(router_wrap_slice_IDATA_4_cfg[31]),
		.out(direct_interc_352_out));

	direct_interc direct_interc_353_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_353_out));

	direct_interc direct_interc_354_ (
		.in(router_wrap_slice_IDATA_4_cfg[32]),
		.out(direct_interc_354_out));

	direct_interc direct_interc_355_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_355_out));

	direct_interc direct_interc_356_ (
		.in(router_wrap_slice_IDATA_4_cfg[33]),
		.out(direct_interc_356_out));

	direct_interc direct_interc_357_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_357_out));

	direct_interc direct_interc_358_ (
		.in(router_wrap_slice_IDATA_4_cfg[34]),
		.out(direct_interc_358_out));

	direct_interc direct_interc_359_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_359_out));

	direct_interc direct_interc_360_ (
		.in(router_wrap_slice_IVALID_0_cfg),
		.out(direct_interc_360_out));

	direct_interc direct_interc_361_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_361_out));

	direct_interc direct_interc_362_ (
		.in(router_wrap_slice_IVALID_1_cfg),
		.out(direct_interc_362_out));

	direct_interc direct_interc_363_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_363_out));

	direct_interc direct_interc_364_ (
		.in(router_wrap_slice_IVALID_2_cfg),
		.out(direct_interc_364_out));

	direct_interc direct_interc_365_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_365_out));

	direct_interc direct_interc_366_ (
		.in(router_wrap_slice_IVALID_3_cfg),
		.out(direct_interc_366_out));

	direct_interc direct_interc_367_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_367_out));

	direct_interc direct_interc_368_ (
		.in(router_wrap_slice_IVALID_4_cfg),
		.out(direct_interc_368_out));

	direct_interc direct_interc_369_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_369_out));

	direct_interc direct_interc_370_ (
		.in(router_wrap_slice_IVCH_0_cfg),
		.out(direct_interc_370_out));

	direct_interc direct_interc_371_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_371_out));

	direct_interc direct_interc_372_ (
		.in(router_wrap_slice_IVCH_1_cfg),
		.out(direct_interc_372_out));

	direct_interc direct_interc_373_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_373_out));

	direct_interc direct_interc_374_ (
		.in(router_wrap_slice_IVCH_2_cfg),
		.out(direct_interc_374_out));

	direct_interc direct_interc_375_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_375_out));

	direct_interc direct_interc_376_ (
		.in(router_wrap_slice_IVCH_3_cfg),
		.out(direct_interc_376_out));

	direct_interc direct_interc_377_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_377_out));

	direct_interc direct_interc_378_ (
		.in(router_wrap_slice_IVCH_4_cfg),
		.out(direct_interc_378_out));

	direct_interc direct_interc_379_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_379_out));

	direct_interc direct_interc_380_ (
		.in(router_wrap_slice_IACK_0_cfg[0]),
		.out(direct_interc_380_out));

	direct_interc direct_interc_381_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_381_out));

	direct_interc direct_interc_382_ (
		.in(router_wrap_slice_IACK_0_cfg[1]),
		.out(direct_interc_382_out));

	direct_interc direct_interc_383_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_383_out));

	direct_interc direct_interc_384_ (
		.in(router_wrap_slice_IACK_1_cfg[0]),
		.out(direct_interc_384_out));

	direct_interc direct_interc_385_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_385_out));

	direct_interc direct_interc_386_ (
		.in(router_wrap_slice_IACK_1_cfg[1]),
		.out(direct_interc_386_out));

	direct_interc direct_interc_387_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_387_out));

	direct_interc direct_interc_388_ (
		.in(router_wrap_slice_IACK_2_cfg[0]),
		.out(direct_interc_388_out));

	direct_interc direct_interc_389_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_389_out));

	direct_interc direct_interc_390_ (
		.in(router_wrap_slice_IACK_2_cfg[1]),
		.out(direct_interc_390_out));

	direct_interc direct_interc_391_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_391_out));

	direct_interc direct_interc_392_ (
		.in(router_wrap_slice_IACK_3_cfg[0]),
		.out(direct_interc_392_out));

	direct_interc direct_interc_393_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_393_out));

	direct_interc direct_interc_394_ (
		.in(router_wrap_slice_IACK_3_cfg[1]),
		.out(direct_interc_394_out));

	direct_interc direct_interc_395_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_395_out));

	direct_interc direct_interc_396_ (
		.in(router_wrap_slice_IACK_4_cfg[0]),
		.out(direct_interc_396_out));

	direct_interc direct_interc_397_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_397_out));

	direct_interc direct_interc_398_ (
		.in(router_wrap_slice_IACK_4_cfg[1]),
		.out(direct_interc_398_out));

	direct_interc direct_interc_399_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_399_out));

	direct_interc direct_interc_400_ (
		.in(router_wrap_slice_ILCK_0_cfg[0]),
		.out(direct_interc_400_out));

	direct_interc direct_interc_401_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_401_out));

	direct_interc direct_interc_402_ (
		.in(router_wrap_slice_ILCK_0_cfg[1]),
		.out(direct_interc_402_out));

	direct_interc direct_interc_403_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_403_out));

	direct_interc direct_interc_404_ (
		.in(router_wrap_slice_ILCK_1_cfg[0]),
		.out(direct_interc_404_out));

	direct_interc direct_interc_405_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_405_out));

	direct_interc direct_interc_406_ (
		.in(router_wrap_slice_ILCK_1_cfg[1]),
		.out(direct_interc_406_out));

	direct_interc direct_interc_407_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_407_out));

	direct_interc direct_interc_408_ (
		.in(router_wrap_slice_ILCK_2_cfg[0]),
		.out(direct_interc_408_out));

	direct_interc direct_interc_409_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_409_out));

	direct_interc direct_interc_410_ (
		.in(router_wrap_slice_ILCK_2_cfg[1]),
		.out(direct_interc_410_out));

	direct_interc direct_interc_411_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_411_out));

	direct_interc direct_interc_412_ (
		.in(router_wrap_slice_ILCK_3_cfg[0]),
		.out(direct_interc_412_out));

	direct_interc direct_interc_413_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_413_out));

	direct_interc direct_interc_414_ (
		.in(router_wrap_slice_ILCK_3_cfg[1]),
		.out(direct_interc_414_out));

	direct_interc direct_interc_415_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_415_out));

	direct_interc direct_interc_416_ (
		.in(router_wrap_slice_ILCK_4_cfg[0]),
		.out(direct_interc_416_out));

	direct_interc direct_interc_417_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_417_out));

	direct_interc direct_interc_418_ (
		.in(router_wrap_slice_ILCK_4_cfg[1]),
		.out(direct_interc_418_out));

	direct_interc direct_interc_419_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_419_out));

	direct_interc direct_interc_420_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[0]),
		.out(direct_interc_420_out));

	direct_interc direct_interc_421_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_421_out));

	direct_interc direct_interc_422_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[1]),
		.out(direct_interc_422_out));

	direct_interc direct_interc_423_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_423_out));

	direct_interc direct_interc_424_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[2]),
		.out(direct_interc_424_out));

	direct_interc direct_interc_425_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_425_out));

	direct_interc direct_interc_426_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[3]),
		.out(direct_interc_426_out));

	direct_interc direct_interc_427_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_427_out));

	direct_interc direct_interc_428_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[4]),
		.out(direct_interc_428_out));

	direct_interc direct_interc_429_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_429_out));

	direct_interc direct_interc_430_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[5]),
		.out(direct_interc_430_out));

	direct_interc direct_interc_431_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_431_out));

	direct_interc direct_interc_432_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[6]),
		.out(direct_interc_432_out));

	direct_interc direct_interc_433_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_433_out));

	direct_interc direct_interc_434_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[7]),
		.out(direct_interc_434_out));

	direct_interc direct_interc_435_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_435_out));

	direct_interc direct_interc_436_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[8]),
		.out(direct_interc_436_out));

	direct_interc direct_interc_437_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_437_out));

	direct_interc direct_interc_438_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[9]),
		.out(direct_interc_438_out));

	direct_interc direct_interc_439_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_439_out));

	direct_interc direct_interc_440_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[10]),
		.out(direct_interc_440_out));

	direct_interc direct_interc_441_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_441_out));

	direct_interc direct_interc_442_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[11]),
		.out(direct_interc_442_out));

	direct_interc direct_interc_443_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_443_out));

	direct_interc direct_interc_444_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[12]),
		.out(direct_interc_444_out));

	direct_interc direct_interc_445_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_445_out));

	direct_interc direct_interc_446_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[13]),
		.out(direct_interc_446_out));

	direct_interc direct_interc_447_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_447_out));

	direct_interc direct_interc_448_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[14]),
		.out(direct_interc_448_out));

	direct_interc direct_interc_449_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_449_out));

	direct_interc direct_interc_450_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[15]),
		.out(direct_interc_450_out));

	direct_interc direct_interc_451_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_451_out));

	direct_interc direct_interc_452_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[16]),
		.out(direct_interc_452_out));

	direct_interc direct_interc_453_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_453_out));

	direct_interc direct_interc_454_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[17]),
		.out(direct_interc_454_out));

	direct_interc direct_interc_455_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_455_out));

	direct_interc direct_interc_456_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[18]),
		.out(direct_interc_456_out));

	direct_interc direct_interc_457_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_457_out));

	direct_interc direct_interc_458_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[19]),
		.out(direct_interc_458_out));

	direct_interc direct_interc_459_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_459_out));

	direct_interc direct_interc_460_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[20]),
		.out(direct_interc_460_out));

	direct_interc direct_interc_461_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_461_out));

	direct_interc direct_interc_462_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[21]),
		.out(direct_interc_462_out));

	direct_interc direct_interc_463_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_463_out));

	direct_interc direct_interc_464_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[22]),
		.out(direct_interc_464_out));

	direct_interc direct_interc_465_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_465_out));

	direct_interc direct_interc_466_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[23]),
		.out(direct_interc_466_out));

	direct_interc direct_interc_467_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_467_out));

	direct_interc direct_interc_468_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[24]),
		.out(direct_interc_468_out));

	direct_interc direct_interc_469_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_469_out));

	direct_interc direct_interc_470_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[25]),
		.out(direct_interc_470_out));

	direct_interc direct_interc_471_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_471_out));

	direct_interc direct_interc_472_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[26]),
		.out(direct_interc_472_out));

	direct_interc direct_interc_473_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_473_out));

	direct_interc direct_interc_474_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[27]),
		.out(direct_interc_474_out));

	direct_interc direct_interc_475_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_475_out));

	direct_interc direct_interc_476_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[28]),
		.out(direct_interc_476_out));

	direct_interc direct_interc_477_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_477_out));

	direct_interc direct_interc_478_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[29]),
		.out(direct_interc_478_out));

	direct_interc direct_interc_479_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_479_out));

	direct_interc direct_interc_480_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[30]),
		.out(direct_interc_480_out));

	direct_interc direct_interc_481_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_481_out));

	direct_interc direct_interc_482_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[31]),
		.out(direct_interc_482_out));

	direct_interc direct_interc_483_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_483_out));

	direct_interc direct_interc_484_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[32]),
		.out(direct_interc_484_out));

	direct_interc direct_interc_485_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_485_out));

	direct_interc direct_interc_486_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[33]),
		.out(direct_interc_486_out));

	direct_interc direct_interc_487_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_487_out));

	direct_interc direct_interc_488_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_0[34]),
		.out(direct_interc_488_out));

	direct_interc direct_interc_489_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_489_out));

	direct_interc direct_interc_490_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[0]),
		.out(direct_interc_490_out));

	direct_interc direct_interc_491_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_491_out));

	direct_interc direct_interc_492_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[1]),
		.out(direct_interc_492_out));

	direct_interc direct_interc_493_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_493_out));

	direct_interc direct_interc_494_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[2]),
		.out(direct_interc_494_out));

	direct_interc direct_interc_495_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_495_out));

	direct_interc direct_interc_496_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[3]),
		.out(direct_interc_496_out));

	direct_interc direct_interc_497_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_497_out));

	direct_interc direct_interc_498_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[4]),
		.out(direct_interc_498_out));

	direct_interc direct_interc_499_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_499_out));

	direct_interc direct_interc_500_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[5]),
		.out(direct_interc_500_out));

	direct_interc direct_interc_501_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_501_out));

	direct_interc direct_interc_502_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[6]),
		.out(direct_interc_502_out));

	direct_interc direct_interc_503_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_503_out));

	direct_interc direct_interc_504_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[7]),
		.out(direct_interc_504_out));

	direct_interc direct_interc_505_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_505_out));

	direct_interc direct_interc_506_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[8]),
		.out(direct_interc_506_out));

	direct_interc direct_interc_507_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_507_out));

	direct_interc direct_interc_508_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[9]),
		.out(direct_interc_508_out));

	direct_interc direct_interc_509_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_509_out));

	direct_interc direct_interc_510_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[10]),
		.out(direct_interc_510_out));

	direct_interc direct_interc_511_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_511_out));

	direct_interc direct_interc_512_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[11]),
		.out(direct_interc_512_out));

	direct_interc direct_interc_513_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_513_out));

	direct_interc direct_interc_514_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[12]),
		.out(direct_interc_514_out));

	direct_interc direct_interc_515_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_515_out));

	direct_interc direct_interc_516_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[13]),
		.out(direct_interc_516_out));

	direct_interc direct_interc_517_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_517_out));

	direct_interc direct_interc_518_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[14]),
		.out(direct_interc_518_out));

	direct_interc direct_interc_519_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_519_out));

	direct_interc direct_interc_520_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[15]),
		.out(direct_interc_520_out));

	direct_interc direct_interc_521_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_521_out));

	direct_interc direct_interc_522_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[16]),
		.out(direct_interc_522_out));

	direct_interc direct_interc_523_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_523_out));

	direct_interc direct_interc_524_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[17]),
		.out(direct_interc_524_out));

	direct_interc direct_interc_525_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_525_out));

	direct_interc direct_interc_526_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[18]),
		.out(direct_interc_526_out));

	direct_interc direct_interc_527_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_527_out));

	direct_interc direct_interc_528_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[19]),
		.out(direct_interc_528_out));

	direct_interc direct_interc_529_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_529_out));

	direct_interc direct_interc_530_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[20]),
		.out(direct_interc_530_out));

	direct_interc direct_interc_531_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_531_out));

	direct_interc direct_interc_532_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[21]),
		.out(direct_interc_532_out));

	direct_interc direct_interc_533_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_533_out));

	direct_interc direct_interc_534_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[22]),
		.out(direct_interc_534_out));

	direct_interc direct_interc_535_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_535_out));

	direct_interc direct_interc_536_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[23]),
		.out(direct_interc_536_out));

	direct_interc direct_interc_537_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_537_out));

	direct_interc direct_interc_538_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[24]),
		.out(direct_interc_538_out));

	direct_interc direct_interc_539_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_539_out));

	direct_interc direct_interc_540_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[25]),
		.out(direct_interc_540_out));

	direct_interc direct_interc_541_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_541_out));

	direct_interc direct_interc_542_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[26]),
		.out(direct_interc_542_out));

	direct_interc direct_interc_543_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_543_out));

	direct_interc direct_interc_544_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[27]),
		.out(direct_interc_544_out));

	direct_interc direct_interc_545_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_545_out));

	direct_interc direct_interc_546_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[28]),
		.out(direct_interc_546_out));

	direct_interc direct_interc_547_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_547_out));

	direct_interc direct_interc_548_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[29]),
		.out(direct_interc_548_out));

	direct_interc direct_interc_549_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_549_out));

	direct_interc direct_interc_550_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[30]),
		.out(direct_interc_550_out));

	direct_interc direct_interc_551_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_551_out));

	direct_interc direct_interc_552_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[31]),
		.out(direct_interc_552_out));

	direct_interc direct_interc_553_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_553_out));

	direct_interc direct_interc_554_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[32]),
		.out(direct_interc_554_out));

	direct_interc direct_interc_555_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_555_out));

	direct_interc direct_interc_556_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[33]),
		.out(direct_interc_556_out));

	direct_interc direct_interc_557_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_557_out));

	direct_interc direct_interc_558_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_1[34]),
		.out(direct_interc_558_out));

	direct_interc direct_interc_559_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_559_out));

	direct_interc direct_interc_560_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[0]),
		.out(direct_interc_560_out));

	direct_interc direct_interc_561_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_561_out));

	direct_interc direct_interc_562_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[1]),
		.out(direct_interc_562_out));

	direct_interc direct_interc_563_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_563_out));

	direct_interc direct_interc_564_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[2]),
		.out(direct_interc_564_out));

	direct_interc direct_interc_565_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_565_out));

	direct_interc direct_interc_566_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[3]),
		.out(direct_interc_566_out));

	direct_interc direct_interc_567_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_567_out));

	direct_interc direct_interc_568_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[4]),
		.out(direct_interc_568_out));

	direct_interc direct_interc_569_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_569_out));

	direct_interc direct_interc_570_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[5]),
		.out(direct_interc_570_out));

	direct_interc direct_interc_571_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_571_out));

	direct_interc direct_interc_572_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[6]),
		.out(direct_interc_572_out));

	direct_interc direct_interc_573_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_573_out));

	direct_interc direct_interc_574_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[7]),
		.out(direct_interc_574_out));

	direct_interc direct_interc_575_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_575_out));

	direct_interc direct_interc_576_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[8]),
		.out(direct_interc_576_out));

	direct_interc direct_interc_577_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_577_out));

	direct_interc direct_interc_578_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[9]),
		.out(direct_interc_578_out));

	direct_interc direct_interc_579_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_579_out));

	direct_interc direct_interc_580_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[10]),
		.out(direct_interc_580_out));

	direct_interc direct_interc_581_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_581_out));

	direct_interc direct_interc_582_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[11]),
		.out(direct_interc_582_out));

	direct_interc direct_interc_583_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_583_out));

	direct_interc direct_interc_584_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[12]),
		.out(direct_interc_584_out));

	direct_interc direct_interc_585_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_585_out));

	direct_interc direct_interc_586_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[13]),
		.out(direct_interc_586_out));

	direct_interc direct_interc_587_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_587_out));

	direct_interc direct_interc_588_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[14]),
		.out(direct_interc_588_out));

	direct_interc direct_interc_589_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_589_out));

	direct_interc direct_interc_590_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[15]),
		.out(direct_interc_590_out));

	direct_interc direct_interc_591_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_591_out));

	direct_interc direct_interc_592_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[16]),
		.out(direct_interc_592_out));

	direct_interc direct_interc_593_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_593_out));

	direct_interc direct_interc_594_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[17]),
		.out(direct_interc_594_out));

	direct_interc direct_interc_595_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_595_out));

	direct_interc direct_interc_596_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[18]),
		.out(direct_interc_596_out));

	direct_interc direct_interc_597_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_597_out));

	direct_interc direct_interc_598_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[19]),
		.out(direct_interc_598_out));

	direct_interc direct_interc_599_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_599_out));

	direct_interc direct_interc_600_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[20]),
		.out(direct_interc_600_out));

	direct_interc direct_interc_601_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_601_out));

	direct_interc direct_interc_602_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[21]),
		.out(direct_interc_602_out));

	direct_interc direct_interc_603_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_603_out));

	direct_interc direct_interc_604_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[22]),
		.out(direct_interc_604_out));

	direct_interc direct_interc_605_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_605_out));

	direct_interc direct_interc_606_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[23]),
		.out(direct_interc_606_out));

	direct_interc direct_interc_607_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_607_out));

	direct_interc direct_interc_608_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[24]),
		.out(direct_interc_608_out));

	direct_interc direct_interc_609_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_609_out));

	direct_interc direct_interc_610_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[25]),
		.out(direct_interc_610_out));

	direct_interc direct_interc_611_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_611_out));

	direct_interc direct_interc_612_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[26]),
		.out(direct_interc_612_out));

	direct_interc direct_interc_613_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_613_out));

	direct_interc direct_interc_614_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[27]),
		.out(direct_interc_614_out));

	direct_interc direct_interc_615_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_615_out));

	direct_interc direct_interc_616_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[28]),
		.out(direct_interc_616_out));

	direct_interc direct_interc_617_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_617_out));

	direct_interc direct_interc_618_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[29]),
		.out(direct_interc_618_out));

	direct_interc direct_interc_619_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_619_out));

	direct_interc direct_interc_620_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[30]),
		.out(direct_interc_620_out));

	direct_interc direct_interc_621_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_621_out));

	direct_interc direct_interc_622_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[31]),
		.out(direct_interc_622_out));

	direct_interc direct_interc_623_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_623_out));

	direct_interc direct_interc_624_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[32]),
		.out(direct_interc_624_out));

	direct_interc direct_interc_625_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_625_out));

	direct_interc direct_interc_626_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[33]),
		.out(direct_interc_626_out));

	direct_interc direct_interc_627_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_627_out));

	direct_interc direct_interc_628_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_2[34]),
		.out(direct_interc_628_out));

	direct_interc direct_interc_629_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_629_out));

	direct_interc direct_interc_630_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[0]),
		.out(direct_interc_630_out));

	direct_interc direct_interc_631_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_631_out));

	direct_interc direct_interc_632_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[1]),
		.out(direct_interc_632_out));

	direct_interc direct_interc_633_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_633_out));

	direct_interc direct_interc_634_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[2]),
		.out(direct_interc_634_out));

	direct_interc direct_interc_635_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_635_out));

	direct_interc direct_interc_636_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[3]),
		.out(direct_interc_636_out));

	direct_interc direct_interc_637_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_637_out));

	direct_interc direct_interc_638_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[4]),
		.out(direct_interc_638_out));

	direct_interc direct_interc_639_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_639_out));

	direct_interc direct_interc_640_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[5]),
		.out(direct_interc_640_out));

	direct_interc direct_interc_641_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_641_out));

	direct_interc direct_interc_642_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[6]),
		.out(direct_interc_642_out));

	direct_interc direct_interc_643_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_643_out));

	direct_interc direct_interc_644_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[7]),
		.out(direct_interc_644_out));

	direct_interc direct_interc_645_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_645_out));

	direct_interc direct_interc_646_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[8]),
		.out(direct_interc_646_out));

	direct_interc direct_interc_647_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_647_out));

	direct_interc direct_interc_648_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[9]),
		.out(direct_interc_648_out));

	direct_interc direct_interc_649_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_649_out));

	direct_interc direct_interc_650_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[10]),
		.out(direct_interc_650_out));

	direct_interc direct_interc_651_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_651_out));

	direct_interc direct_interc_652_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[11]),
		.out(direct_interc_652_out));

	direct_interc direct_interc_653_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_653_out));

	direct_interc direct_interc_654_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[12]),
		.out(direct_interc_654_out));

	direct_interc direct_interc_655_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_655_out));

	direct_interc direct_interc_656_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[13]),
		.out(direct_interc_656_out));

	direct_interc direct_interc_657_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_657_out));

	direct_interc direct_interc_658_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[14]),
		.out(direct_interc_658_out));

	direct_interc direct_interc_659_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_659_out));

	direct_interc direct_interc_660_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[15]),
		.out(direct_interc_660_out));

	direct_interc direct_interc_661_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_661_out));

	direct_interc direct_interc_662_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[16]),
		.out(direct_interc_662_out));

	direct_interc direct_interc_663_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_663_out));

	direct_interc direct_interc_664_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[17]),
		.out(direct_interc_664_out));

	direct_interc direct_interc_665_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_665_out));

	direct_interc direct_interc_666_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[18]),
		.out(direct_interc_666_out));

	direct_interc direct_interc_667_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_667_out));

	direct_interc direct_interc_668_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[19]),
		.out(direct_interc_668_out));

	direct_interc direct_interc_669_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_669_out));

	direct_interc direct_interc_670_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[20]),
		.out(direct_interc_670_out));

	direct_interc direct_interc_671_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_671_out));

	direct_interc direct_interc_672_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[21]),
		.out(direct_interc_672_out));

	direct_interc direct_interc_673_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_673_out));

	direct_interc direct_interc_674_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[22]),
		.out(direct_interc_674_out));

	direct_interc direct_interc_675_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_675_out));

	direct_interc direct_interc_676_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[23]),
		.out(direct_interc_676_out));

	direct_interc direct_interc_677_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_677_out));

	direct_interc direct_interc_678_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[24]),
		.out(direct_interc_678_out));

	direct_interc direct_interc_679_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_679_out));

	direct_interc direct_interc_680_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[25]),
		.out(direct_interc_680_out));

	direct_interc direct_interc_681_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_681_out));

	direct_interc direct_interc_682_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[26]),
		.out(direct_interc_682_out));

	direct_interc direct_interc_683_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_683_out));

	direct_interc direct_interc_684_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[27]),
		.out(direct_interc_684_out));

	direct_interc direct_interc_685_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_685_out));

	direct_interc direct_interc_686_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[28]),
		.out(direct_interc_686_out));

	direct_interc direct_interc_687_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_687_out));

	direct_interc direct_interc_688_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[29]),
		.out(direct_interc_688_out));

	direct_interc direct_interc_689_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_689_out));

	direct_interc direct_interc_690_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[30]),
		.out(direct_interc_690_out));

	direct_interc direct_interc_691_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_691_out));

	direct_interc direct_interc_692_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[31]),
		.out(direct_interc_692_out));

	direct_interc direct_interc_693_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_693_out));

	direct_interc direct_interc_694_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[32]),
		.out(direct_interc_694_out));

	direct_interc direct_interc_695_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_695_out));

	direct_interc direct_interc_696_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[33]),
		.out(direct_interc_696_out));

	direct_interc direct_interc_697_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_697_out));

	direct_interc direct_interc_698_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_3[34]),
		.out(direct_interc_698_out));

	direct_interc direct_interc_699_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_699_out));

	direct_interc direct_interc_700_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[0]),
		.out(direct_interc_700_out));

	direct_interc direct_interc_701_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_701_out));

	direct_interc direct_interc_702_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[1]),
		.out(direct_interc_702_out));

	direct_interc direct_interc_703_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_703_out));

	direct_interc direct_interc_704_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[2]),
		.out(direct_interc_704_out));

	direct_interc direct_interc_705_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_705_out));

	direct_interc direct_interc_706_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[3]),
		.out(direct_interc_706_out));

	direct_interc direct_interc_707_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_707_out));

	direct_interc direct_interc_708_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[4]),
		.out(direct_interc_708_out));

	direct_interc direct_interc_709_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_709_out));

	direct_interc direct_interc_710_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[5]),
		.out(direct_interc_710_out));

	direct_interc direct_interc_711_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_711_out));

	direct_interc direct_interc_712_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[6]),
		.out(direct_interc_712_out));

	direct_interc direct_interc_713_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_713_out));

	direct_interc direct_interc_714_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[7]),
		.out(direct_interc_714_out));

	direct_interc direct_interc_715_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_715_out));

	direct_interc direct_interc_716_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[8]),
		.out(direct_interc_716_out));

	direct_interc direct_interc_717_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_717_out));

	direct_interc direct_interc_718_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[9]),
		.out(direct_interc_718_out));

	direct_interc direct_interc_719_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_719_out));

	direct_interc direct_interc_720_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[10]),
		.out(direct_interc_720_out));

	direct_interc direct_interc_721_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_721_out));

	direct_interc direct_interc_722_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[11]),
		.out(direct_interc_722_out));

	direct_interc direct_interc_723_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_723_out));

	direct_interc direct_interc_724_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[12]),
		.out(direct_interc_724_out));

	direct_interc direct_interc_725_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_725_out));

	direct_interc direct_interc_726_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[13]),
		.out(direct_interc_726_out));

	direct_interc direct_interc_727_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_727_out));

	direct_interc direct_interc_728_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[14]),
		.out(direct_interc_728_out));

	direct_interc direct_interc_729_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_729_out));

	direct_interc direct_interc_730_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[15]),
		.out(direct_interc_730_out));

	direct_interc direct_interc_731_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_731_out));

	direct_interc direct_interc_732_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[16]),
		.out(direct_interc_732_out));

	direct_interc direct_interc_733_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_733_out));

	direct_interc direct_interc_734_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[17]),
		.out(direct_interc_734_out));

	direct_interc direct_interc_735_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_735_out));

	direct_interc direct_interc_736_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[18]),
		.out(direct_interc_736_out));

	direct_interc direct_interc_737_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_737_out));

	direct_interc direct_interc_738_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[19]),
		.out(direct_interc_738_out));

	direct_interc direct_interc_739_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_739_out));

	direct_interc direct_interc_740_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[20]),
		.out(direct_interc_740_out));

	direct_interc direct_interc_741_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_741_out));

	direct_interc direct_interc_742_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[21]),
		.out(direct_interc_742_out));

	direct_interc direct_interc_743_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_743_out));

	direct_interc direct_interc_744_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[22]),
		.out(direct_interc_744_out));

	direct_interc direct_interc_745_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_745_out));

	direct_interc direct_interc_746_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[23]),
		.out(direct_interc_746_out));

	direct_interc direct_interc_747_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_747_out));

	direct_interc direct_interc_748_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[24]),
		.out(direct_interc_748_out));

	direct_interc direct_interc_749_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_749_out));

	direct_interc direct_interc_750_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[25]),
		.out(direct_interc_750_out));

	direct_interc direct_interc_751_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_751_out));

	direct_interc direct_interc_752_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[26]),
		.out(direct_interc_752_out));

	direct_interc direct_interc_753_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_753_out));

	direct_interc direct_interc_754_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[27]),
		.out(direct_interc_754_out));

	direct_interc direct_interc_755_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_755_out));

	direct_interc direct_interc_756_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[28]),
		.out(direct_interc_756_out));

	direct_interc direct_interc_757_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_757_out));

	direct_interc direct_interc_758_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[29]),
		.out(direct_interc_758_out));

	direct_interc direct_interc_759_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_759_out));

	direct_interc direct_interc_760_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[30]),
		.out(direct_interc_760_out));

	direct_interc direct_interc_761_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_761_out));

	direct_interc direct_interc_762_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[31]),
		.out(direct_interc_762_out));

	direct_interc direct_interc_763_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_763_out));

	direct_interc direct_interc_764_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[32]),
		.out(direct_interc_764_out));

	direct_interc direct_interc_765_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_765_out));

	direct_interc direct_interc_766_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[33]),
		.out(direct_interc_766_out));

	direct_interc direct_interc_767_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_767_out));

	direct_interc direct_interc_768_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ODATA_4[34]),
		.out(direct_interc_768_out));

	direct_interc direct_interc_769_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_769_out));

	direct_interc direct_interc_770_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_0),
		.out(direct_interc_770_out));

	direct_interc direct_interc_771_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_771_out));

	direct_interc direct_interc_772_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_1),
		.out(direct_interc_772_out));

	direct_interc direct_interc_773_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_773_out));

	direct_interc direct_interc_774_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_2),
		.out(direct_interc_774_out));

	direct_interc direct_interc_775_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_775_out));

	direct_interc direct_interc_776_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_3),
		.out(direct_interc_776_out));

	direct_interc direct_interc_777_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_777_out));

	direct_interc direct_interc_778_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVALID_4),
		.out(direct_interc_778_out));

	direct_interc direct_interc_779_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_779_out));

	direct_interc direct_interc_780_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_0),
		.out(direct_interc_780_out));

	direct_interc direct_interc_781_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_781_out));

	direct_interc direct_interc_782_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_1),
		.out(direct_interc_782_out));

	direct_interc direct_interc_783_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_783_out));

	direct_interc direct_interc_784_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_2),
		.out(direct_interc_784_out));

	direct_interc direct_interc_785_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_785_out));

	direct_interc direct_interc_786_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_3),
		.out(direct_interc_786_out));

	direct_interc direct_interc_787_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_787_out));

	direct_interc direct_interc_788_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OVCH_4),
		.out(direct_interc_788_out));

	direct_interc direct_interc_789_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_789_out));

	direct_interc direct_interc_790_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0[0]),
		.out(direct_interc_790_out));

	direct_interc direct_interc_791_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_791_out));

	direct_interc direct_interc_792_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_0[1]),
		.out(direct_interc_792_out));

	direct_interc direct_interc_793_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_793_out));

	direct_interc direct_interc_794_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1[0]),
		.out(direct_interc_794_out));

	direct_interc direct_interc_795_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_795_out));

	direct_interc direct_interc_796_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_1[1]),
		.out(direct_interc_796_out));

	direct_interc direct_interc_797_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_797_out));

	direct_interc direct_interc_798_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2[0]),
		.out(direct_interc_798_out));

	direct_interc direct_interc_799_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_799_out));

	direct_interc direct_interc_800_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_2[1]),
		.out(direct_interc_800_out));

	direct_interc direct_interc_801_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_801_out));

	direct_interc direct_interc_802_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3[0]),
		.out(direct_interc_802_out));

	direct_interc direct_interc_803_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_803_out));

	direct_interc direct_interc_804_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_3[1]),
		.out(direct_interc_804_out));

	direct_interc direct_interc_805_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_805_out));

	direct_interc direct_interc_806_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4[0]),
		.out(direct_interc_806_out));

	direct_interc direct_interc_807_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_807_out));

	direct_interc direct_interc_808_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OACK_4[1]),
		.out(direct_interc_808_out));

	direct_interc direct_interc_809_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_809_out));

	direct_interc direct_interc_810_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0[0]),
		.out(direct_interc_810_out));

	direct_interc direct_interc_811_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_811_out));

	direct_interc direct_interc_812_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_0[1]),
		.out(direct_interc_812_out));

	direct_interc direct_interc_813_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_813_out));

	direct_interc direct_interc_814_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1[0]),
		.out(direct_interc_814_out));

	direct_interc direct_interc_815_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_815_out));

	direct_interc direct_interc_816_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_1[1]),
		.out(direct_interc_816_out));

	direct_interc direct_interc_817_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_817_out));

	direct_interc direct_interc_818_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2[0]),
		.out(direct_interc_818_out));

	direct_interc direct_interc_819_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_819_out));

	direct_interc direct_interc_820_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_2[1]),
		.out(direct_interc_820_out));

	direct_interc direct_interc_821_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_821_out));

	direct_interc direct_interc_822_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3[0]),
		.out(direct_interc_822_out));

	direct_interc direct_interc_823_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_823_out));

	direct_interc direct_interc_824_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_3[1]),
		.out(direct_interc_824_out));

	direct_interc direct_interc_825_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_825_out));

	direct_interc direct_interc_826_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4[0]),
		.out(direct_interc_826_out));

	direct_interc direct_interc_827_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_827_out));

	direct_interc direct_interc_828_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_ORDY_4[1]),
		.out(direct_interc_828_out));

	direct_interc direct_interc_829_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_829_out));

	direct_interc direct_interc_830_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0[0]),
		.out(direct_interc_830_out));

	direct_interc direct_interc_831_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_831_out));

	direct_interc direct_interc_832_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_0[1]),
		.out(direct_interc_832_out));

	direct_interc direct_interc_833_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_833_out));

	direct_interc direct_interc_834_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1[0]),
		.out(direct_interc_834_out));

	direct_interc direct_interc_835_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_835_out));

	direct_interc direct_interc_836_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_1[1]),
		.out(direct_interc_836_out));

	direct_interc direct_interc_837_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_837_out));

	direct_interc direct_interc_838_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2[0]),
		.out(direct_interc_838_out));

	direct_interc direct_interc_839_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_839_out));

	direct_interc direct_interc_840_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_2[1]),
		.out(direct_interc_840_out));

	direct_interc direct_interc_841_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_841_out));

	direct_interc direct_interc_842_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3[0]),
		.out(direct_interc_842_out));

	direct_interc direct_interc_843_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_843_out));

	direct_interc direct_interc_844_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_3[1]),
		.out(direct_interc_844_out));

	direct_interc direct_interc_845_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_845_out));

	direct_interc direct_interc_846_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4[0]),
		.out(direct_interc_846_out));

	direct_interc direct_interc_847_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_847_out));

	direct_interc direct_interc_848_ (
		.in(logical_tile_router_mode_router_wrap__router_wrap_slice_mode_default__router_wrap_0_router_wrap_OLCK_4[1]),
		.out(direct_interc_848_out));

	direct_interc direct_interc_849_ (
		.in(router_wrap_slice_clk),
		.out(direct_interc_849_out));

endmodule
// ----- END Verilog module for logical_tile_router_mode_router_wrap__router_wrap_slice -----

//----- Default net type -----
`default_nettype wire



// ----- END Physical programmable logic block Verilog module: router_wrap_slice -----
