//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[18][16]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Jul 20 12:17:04 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_18__16_ -----
module sb_18__16_(prog_clk,
                  chany_top_in,
                  top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                  top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                  top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                  chany_bottom_in,
                  bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                  bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                  bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_,
                  chanx_left_in,
                  left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                  left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                  left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                  ccff_head,
                  chany_top_out,
                  chany_bottom_out,
                  chanx_left_out,
                  ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:160] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:160] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_;
//----- INPUT PORTS -----
input [0:160] chanx_left_in;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:160] chany_top_out;
//----- OUTPUT PORTS -----
output [0:160] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:160] chanx_left_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_100_sram;
wire [0:1] mux_tree_tapbuf_size3_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_101_sram;
wire [0:1] mux_tree_tapbuf_size3_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_102_sram;
wire [0:1] mux_tree_tapbuf_size3_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_103_sram;
wire [0:1] mux_tree_tapbuf_size3_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_104_sram;
wire [0:1] mux_tree_tapbuf_size3_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_105_sram;
wire [0:1] mux_tree_tapbuf_size3_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_106_sram;
wire [0:1] mux_tree_tapbuf_size3_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_107_sram;
wire [0:1] mux_tree_tapbuf_size3_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_108_sram;
wire [0:1] mux_tree_tapbuf_size3_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_109_sram;
wire [0:1] mux_tree_tapbuf_size3_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_110_sram;
wire [0:1] mux_tree_tapbuf_size3_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_111_sram;
wire [0:1] mux_tree_tapbuf_size3_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_112_sram;
wire [0:1] mux_tree_tapbuf_size3_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_113_sram;
wire [0:1] mux_tree_tapbuf_size3_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_114_sram;
wire [0:1] mux_tree_tapbuf_size3_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_115_sram;
wire [0:1] mux_tree_tapbuf_size3_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_116_sram;
wire [0:1] mux_tree_tapbuf_size3_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_117_sram;
wire [0:1] mux_tree_tapbuf_size3_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_118_sram;
wire [0:1] mux_tree_tapbuf_size3_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_119_sram;
wire [0:1] mux_tree_tapbuf_size3_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_120_sram;
wire [0:1] mux_tree_tapbuf_size3_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_121_sram;
wire [0:1] mux_tree_tapbuf_size3_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_122_sram;
wire [0:1] mux_tree_tapbuf_size3_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_123_sram;
wire [0:1] mux_tree_tapbuf_size3_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_124_sram;
wire [0:1] mux_tree_tapbuf_size3_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_125_sram;
wire [0:1] mux_tree_tapbuf_size3_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_126_sram;
wire [0:1] mux_tree_tapbuf_size3_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_127_sram;
wire [0:1] mux_tree_tapbuf_size3_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_128_sram;
wire [0:1] mux_tree_tapbuf_size3_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_129_sram;
wire [0:1] mux_tree_tapbuf_size3_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_130_sram;
wire [0:1] mux_tree_tapbuf_size3_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_131_sram;
wire [0:1] mux_tree_tapbuf_size3_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_132_sram;
wire [0:1] mux_tree_tapbuf_size3_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_133_sram;
wire [0:1] mux_tree_tapbuf_size3_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_134_sram;
wire [0:1] mux_tree_tapbuf_size3_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_135_sram;
wire [0:1] mux_tree_tapbuf_size3_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_136_sram;
wire [0:1] mux_tree_tapbuf_size3_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_60_sram;
wire [0:1] mux_tree_tapbuf_size3_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_61_sram;
wire [0:1] mux_tree_tapbuf_size3_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_62_sram;
wire [0:1] mux_tree_tapbuf_size3_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_63_sram;
wire [0:1] mux_tree_tapbuf_size3_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_64_sram;
wire [0:1] mux_tree_tapbuf_size3_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_65_sram;
wire [0:1] mux_tree_tapbuf_size3_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_66_sram;
wire [0:1] mux_tree_tapbuf_size3_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_67_sram;
wire [0:1] mux_tree_tapbuf_size3_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_68_sram;
wire [0:1] mux_tree_tapbuf_size3_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_69_sram;
wire [0:1] mux_tree_tapbuf_size3_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_70_sram;
wire [0:1] mux_tree_tapbuf_size3_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_71_sram;
wire [0:1] mux_tree_tapbuf_size3_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_72_sram;
wire [0:1] mux_tree_tapbuf_size3_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_73_sram;
wire [0:1] mux_tree_tapbuf_size3_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_74_sram;
wire [0:1] mux_tree_tapbuf_size3_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_75_sram;
wire [0:1] mux_tree_tapbuf_size3_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_76_sram;
wire [0:1] mux_tree_tapbuf_size3_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_77_sram;
wire [0:1] mux_tree_tapbuf_size3_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_78_sram;
wire [0:1] mux_tree_tapbuf_size3_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_79_sram;
wire [0:1] mux_tree_tapbuf_size3_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_80_sram;
wire [0:1] mux_tree_tapbuf_size3_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_81_sram;
wire [0:1] mux_tree_tapbuf_size3_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_82_sram;
wire [0:1] mux_tree_tapbuf_size3_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_83_sram;
wire [0:1] mux_tree_tapbuf_size3_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_84_sram;
wire [0:1] mux_tree_tapbuf_size3_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_85_sram;
wire [0:1] mux_tree_tapbuf_size3_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_86_sram;
wire [0:1] mux_tree_tapbuf_size3_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_87_sram;
wire [0:1] mux_tree_tapbuf_size3_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_88_sram;
wire [0:1] mux_tree_tapbuf_size3_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_89_sram;
wire [0:1] mux_tree_tapbuf_size3_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_90_sram;
wire [0:1] mux_tree_tapbuf_size3_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_91_sram;
wire [0:1] mux_tree_tapbuf_size3_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_92_sram;
wire [0:1] mux_tree_tapbuf_size3_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_93_sram;
wire [0:1] mux_tree_tapbuf_size3_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_94_sram;
wire [0:1] mux_tree_tapbuf_size3_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_95_sram;
wire [0:1] mux_tree_tapbuf_size3_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_96_sram;
wire [0:1] mux_tree_tapbuf_size3_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_97_sram;
wire [0:1] mux_tree_tapbuf_size3_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_98_sram;
wire [0:1] mux_tree_tapbuf_size3_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_99_sram;
wire [0:1] mux_tree_tapbuf_size3_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_10_sram;
wire [0:2] mux_tree_tapbuf_size4_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_4_sram;
wire [0:2] mux_tree_tapbuf_size4_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_5_sram;
wire [0:2] mux_tree_tapbuf_size4_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_6_sram;
wire [0:2] mux_tree_tapbuf_size4_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_7_sram;
wire [0:2] mux_tree_tapbuf_size4_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_8_sram;
wire [0:2] mux_tree_tapbuf_size4_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_9_sram;
wire [0:2] mux_tree_tapbuf_size4_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_10_sram;
wire [0:2] mux_tree_tapbuf_size5_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_11_sram;
wire [0:2] mux_tree_tapbuf_size5_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_12_sram;
wire [0:2] mux_tree_tapbuf_size5_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_13_sram;
wire [0:2] mux_tree_tapbuf_size5_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_14_sram;
wire [0:2] mux_tree_tapbuf_size5_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_15_sram;
wire [0:2] mux_tree_tapbuf_size5_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_16_sram;
wire [0:2] mux_tree_tapbuf_size5_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_17_sram;
wire [0:2] mux_tree_tapbuf_size5_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_18_sram;
wire [0:2] mux_tree_tapbuf_size5_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_19_sram;
wire [0:2] mux_tree_tapbuf_size5_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_20_sram;
wire [0:2] mux_tree_tapbuf_size5_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_21_sram;
wire [0:2] mux_tree_tapbuf_size5_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_22_sram;
wire [0:2] mux_tree_tapbuf_size5_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_23_sram;
wire [0:2] mux_tree_tapbuf_size5_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_24_sram;
wire [0:2] mux_tree_tapbuf_size5_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_7_sram;
wire [0:2] mux_tree_tapbuf_size5_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_8_sram;
wire [0:2] mux_tree_tapbuf_size5_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_9_sram;
wire [0:2] mux_tree_tapbuf_size5_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_11_sram;
wire [0:2] mux_tree_tapbuf_size6_11_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_12_sram;
wire [0:2] mux_tree_tapbuf_size6_12_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_13_sram;
wire [0:2] mux_tree_tapbuf_size6_13_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_14_sram;
wire [0:2] mux_tree_tapbuf_size6_14_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_15_sram;
wire [0:2] mux_tree_tapbuf_size6_15_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_16_sram;
wire [0:2] mux_tree_tapbuf_size6_16_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_17_sram;
wire [0:2] mux_tree_tapbuf_size6_17_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_18_sram;
wire [0:2] mux_tree_tapbuf_size6_18_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_19_sram;
wire [0:2] mux_tree_tapbuf_size6_19_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_20_sram;
wire [0:2] mux_tree_tapbuf_size6_20_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_21_sram;
wire [0:2] mux_tree_tapbuf_size6_21_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_22_sram;
wire [0:2] mux_tree_tapbuf_size6_22_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_23_sram;
wire [0:2] mux_tree_tapbuf_size6_23_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_24_sram;
wire [0:2] mux_tree_tapbuf_size6_24_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_25_sram;
wire [0:2] mux_tree_tapbuf_size6_25_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_26_sram;
wire [0:2] mux_tree_tapbuf_size6_26_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_27_sram;
wire [0:2] mux_tree_tapbuf_size6_27_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_28_sram;
wire [0:2] mux_tree_tapbuf_size6_28_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_29_sram;
wire [0:2] mux_tree_tapbuf_size6_29_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_30_sram;
wire [0:2] mux_tree_tapbuf_size6_30_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_31_sram;
wire [0:2] mux_tree_tapbuf_size6_31_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_32_sram;
wire [0:2] mux_tree_tapbuf_size6_32_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_33_sram;
wire [0:2] mux_tree_tapbuf_size6_33_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_34_sram;
wire [0:2] mux_tree_tapbuf_size6_34_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_35_sram;
wire [0:2] mux_tree_tapbuf_size6_35_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_36_sram;
wire [0:2] mux_tree_tapbuf_size6_36_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_37_sram;
wire [0:2] mux_tree_tapbuf_size6_37_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_38_sram;
wire [0:2] mux_tree_tapbuf_size6_38_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_39_sram;
wire [0:2] mux_tree_tapbuf_size6_39_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_40_sram;
wire [0:2] mux_tree_tapbuf_size6_40_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_41_sram;
wire [0:2] mux_tree_tapbuf_size6_41_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_42_sram;
wire [0:2] mux_tree_tapbuf_size6_42_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_10_sram;
wire [0:2] mux_tree_tapbuf_size7_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_3_sram;
wire [0:2] mux_tree_tapbuf_size7_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_4_sram;
wire [0:2] mux_tree_tapbuf_size7_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_5_sram;
wire [0:2] mux_tree_tapbuf_size7_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_6_sram;
wire [0:2] mux_tree_tapbuf_size7_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_7_sram;
wire [0:2] mux_tree_tapbuf_size7_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_8_sram;
wire [0:2] mux_tree_tapbuf_size7_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_9_sram;
wire [0:2] mux_tree_tapbuf_size7_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_9_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 72 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[73] = chany_top_in[72];
// ----- Local connection due to Wire 73 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[74] = chany_top_in[73];
// ----- Local connection due to Wire 74 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[75] = chany_top_in[74];
// ----- Local connection due to Wire 76 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[77] = chany_top_in[76];
// ----- Local connection due to Wire 77 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[78] = chany_top_in[77];
// ----- Local connection due to Wire 78 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[79] = chany_top_in[78];
// ----- Local connection due to Wire 80 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[81] = chany_top_in[80];
// ----- Local connection due to Wire 81 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[82] = chany_top_in[81];
// ----- Local connection due to Wire 82 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[83] = chany_top_in[82];
// ----- Local connection due to Wire 84 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[85] = chany_top_in[84];
// ----- Local connection due to Wire 85 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[86] = chany_top_in[85];
// ----- Local connection due to Wire 86 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[87] = chany_top_in[86];
// ----- Local connection due to Wire 88 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[89] = chany_top_in[88];
// ----- Local connection due to Wire 89 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[90] = chany_top_in[89];
// ----- Local connection due to Wire 90 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[91] = chany_top_in[90];
// ----- Local connection due to Wire 92 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[93] = chany_top_in[92];
// ----- Local connection due to Wire 93 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[94] = chany_top_in[93];
// ----- Local connection due to Wire 94 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[95] = chany_top_in[94];
// ----- Local connection due to Wire 96 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[97] = chany_top_in[96];
// ----- Local connection due to Wire 97 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[98] = chany_top_in[97];
// ----- Local connection due to Wire 98 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[99] = chany_top_in[98];
// ----- Local connection due to Wire 100 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[101] = chany_top_in[100];
// ----- Local connection due to Wire 101 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[102] = chany_top_in[101];
// ----- Local connection due to Wire 102 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[103] = chany_top_in[102];
// ----- Local connection due to Wire 104 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[105] = chany_top_in[104];
// ----- Local connection due to Wire 105 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[106] = chany_top_in[105];
// ----- Local connection due to Wire 106 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[107] = chany_top_in[106];
// ----- Local connection due to Wire 108 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[109] = chany_top_in[108];
// ----- Local connection due to Wire 109 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[110] = chany_top_in[109];
// ----- Local connection due to Wire 110 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[111] = chany_top_in[110];
// ----- Local connection due to Wire 112 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[113] = chany_top_in[112];
// ----- Local connection due to Wire 113 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[114] = chany_top_in[113];
// ----- Local connection due to Wire 114 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[115] = chany_top_in[114];
// ----- Local connection due to Wire 116 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[117] = chany_top_in[116];
// ----- Local connection due to Wire 117 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[118] = chany_top_in[117];
// ----- Local connection due to Wire 118 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[119] = chany_top_in[118];
// ----- Local connection due to Wire 120 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[121] = chany_top_in[120];
// ----- Local connection due to Wire 121 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[122] = chany_top_in[121];
// ----- Local connection due to Wire 122 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[123] = chany_top_in[122];
// ----- Local connection due to Wire 124 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[125] = chany_top_in[124];
// ----- Local connection due to Wire 125 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[126] = chany_top_in[125];
// ----- Local connection due to Wire 126 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[127] = chany_top_in[126];
// ----- Local connection due to Wire 128 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[129] = chany_top_in[128];
// ----- Local connection due to Wire 129 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[130] = chany_top_in[129];
// ----- Local connection due to Wire 130 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[131] = chany_top_in[130];
// ----- Local connection due to Wire 132 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[133] = chany_top_in[132];
// ----- Local connection due to Wire 133 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[134] = chany_top_in[133];
// ----- Local connection due to Wire 134 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[135] = chany_top_in[134];
// ----- Local connection due to Wire 136 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[137] = chany_top_in[136];
// ----- Local connection due to Wire 137 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[138] = chany_top_in[137];
// ----- Local connection due to Wire 138 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[139] = chany_top_in[138];
// ----- Local connection due to Wire 140 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[141] = chany_top_in[140];
// ----- Local connection due to Wire 141 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[142] = chany_top_in[141];
// ----- Local connection due to Wire 142 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[143] = chany_top_in[142];
// ----- Local connection due to Wire 144 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[145] = chany_top_in[144];
// ----- Local connection due to Wire 145 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[146] = chany_top_in[145];
// ----- Local connection due to Wire 146 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[147] = chany_top_in[146];
// ----- Local connection due to Wire 148 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[149] = chany_top_in[148];
// ----- Local connection due to Wire 149 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[150] = chany_top_in[149];
// ----- Local connection due to Wire 150 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[151] = chany_top_in[150];
// ----- Local connection due to Wire 152 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[153] = chany_top_in[152];
// ----- Local connection due to Wire 153 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[154] = chany_top_in[153];
// ----- Local connection due to Wire 154 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[155] = chany_top_in[154];
// ----- Local connection due to Wire 156 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[157] = chany_top_in[156];
// ----- Local connection due to Wire 157 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[158] = chany_top_in[157];
// ----- Local connection due to Wire 158 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_bottom_out[159] = chany_top_in[158];
// ----- Local connection due to Wire 177 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 178 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 179 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 181 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 182 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 183 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 185 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 186 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 187 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 189 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 190 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 191 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 193 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 194 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 195 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 197 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 198 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 199 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 201 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 202 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 203 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 205 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 206 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 207 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 209 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 210 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 211 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 213 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 214 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 215 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 217 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 218 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 219 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 221 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 222 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 223 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 225 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 226 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 227 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 229 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 230 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 231 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 233 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 234 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 235 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 237 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 238 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 239 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 241 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 242 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 246 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[73] = chany_bottom_in[72];
// ----- Local connection due to Wire 250 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[74] = chany_bottom_in[73];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[75] = chany_bottom_in[74];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[77] = chany_bottom_in[76];
// ----- Local connection due to Wire 254 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[78] = chany_bottom_in[77];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[79] = chany_bottom_in[78];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[81] = chany_bottom_in[80];
// ----- Local connection due to Wire 258 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[82] = chany_bottom_in[81];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[83] = chany_bottom_in[82];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[85] = chany_bottom_in[84];
// ----- Local connection due to Wire 262 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[86] = chany_bottom_in[85];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[87] = chany_bottom_in[86];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[89] = chany_bottom_in[88];
// ----- Local connection due to Wire 266 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[90] = chany_bottom_in[89];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[91] = chany_bottom_in[90];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[93] = chany_bottom_in[92];
// ----- Local connection due to Wire 270 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[94] = chany_bottom_in[93];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[95] = chany_bottom_in[94];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[97] = chany_bottom_in[96];
// ----- Local connection due to Wire 274 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[98] = chany_bottom_in[97];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[99] = chany_bottom_in[98];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[101] = chany_bottom_in[100];
// ----- Local connection due to Wire 278 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[102] = chany_bottom_in[101];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[103] = chany_bottom_in[102];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[105] = chany_bottom_in[104];
// ----- Local connection due to Wire 282 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[106] = chany_bottom_in[105];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[107] = chany_bottom_in[106];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[109] = chany_bottom_in[108];
// ----- Local connection due to Wire 286 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[110] = chany_bottom_in[109];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[111] = chany_bottom_in[110];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[113] = chany_bottom_in[112];
// ----- Local connection due to Wire 290 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[114] = chany_bottom_in[113];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[115] = chany_bottom_in[114];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[117] = chany_bottom_in[116];
// ----- Local connection due to Wire 294 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[118] = chany_bottom_in[117];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[119] = chany_bottom_in[118];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[121] = chany_bottom_in[120];
// ----- Local connection due to Wire 298 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[122] = chany_bottom_in[121];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[123] = chany_bottom_in[122];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[125] = chany_bottom_in[124];
// ----- Local connection due to Wire 302 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[126] = chany_bottom_in[125];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[127] = chany_bottom_in[126];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[129] = chany_bottom_in[128];
// ----- Local connection due to Wire 306 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[130] = chany_bottom_in[129];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[131] = chany_bottom_in[130];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[133] = chany_bottom_in[132];
// ----- Local connection due to Wire 310 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[134] = chany_bottom_in[133];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[135] = chany_bottom_in[134];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[137] = chany_bottom_in[136];
// ----- Local connection due to Wire 314 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[138] = chany_bottom_in[137];
// ----- Local connection due to Wire 315 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[139] = chany_bottom_in[138];
// ----- Local connection due to Wire 317 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[141] = chany_bottom_in[140];
// ----- Local connection due to Wire 318 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[142] = chany_bottom_in[141];
// ----- Local connection due to Wire 319 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[143] = chany_bottom_in[142];
// ----- Local connection due to Wire 321 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[145] = chany_bottom_in[144];
// ----- Local connection due to Wire 322 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[146] = chany_bottom_in[145];
// ----- Local connection due to Wire 323 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[147] = chany_bottom_in[146];
// ----- Local connection due to Wire 325 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[149] = chany_bottom_in[148];
// ----- Local connection due to Wire 326 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[150] = chany_bottom_in[149];
// ----- Local connection due to Wire 327 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[151] = chany_bottom_in[150];
// ----- Local connection due to Wire 329 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[153] = chany_bottom_in[152];
// ----- Local connection due to Wire 330 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[154] = chany_bottom_in[153];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[155] = chany_bottom_in[154];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[157] = chany_bottom_in[156];
// ----- Local connection due to Wire 334 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[158] = chany_bottom_in[157];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[159] = chany_bottom_in[158];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size7 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[0], chanx_left_in[41], chanx_left_in[82], chanx_left_in[123]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size7 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[37], chanx_left_in[78], chanx_left_in[119], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size7 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[36], chanx_left_in[77], chanx_left_in[118], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size7 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[35], chanx_left_in[76], chanx_left_in[117], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size7_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_3_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size7 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[33], chanx_left_in[74], chanx_left_in[115], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size7_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_4_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size7 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[32], chanx_left_in[73], chanx_left_in[114], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size7_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_5_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size7 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[31], chanx_left_in[72], chanx_left_in[113], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size7_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_6_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size7 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[30], chanx_left_in[71], chanx_left_in[112], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size7_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_7_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size7 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[29], chanx_left_in[70], chanx_left_in[111], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size7_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_8_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size7 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[28], chanx_left_in[69], chanx_left_in[110], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size7_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_9_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size7 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[27], chanx_left_in[68], chanx_left_in[109], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size7_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_10_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size7_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_3_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_4_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_5_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_6_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_7_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_8_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_9_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_10_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[40], chanx_left_in[81], chanx_left_in[122]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size6 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[39], chanx_left_in[80], chanx_left_in[121]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size6 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[38], chanx_left_in[79], chanx_left_in[120]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size6 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[34], chanx_left_in[75], chanx_left_in[116], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size6 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[26], chanx_left_in[67], chanx_left_in[108], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size6 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[25], chanx_left_in[66], chanx_left_in[107], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size6 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[24], chanx_left_in[65], chanx_left_in[106], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[23], chanx_left_in[64], chanx_left_in[105], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size6 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[22], chanx_left_in[63], chanx_left_in[104], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size6 mux_top_track_160 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[21], chanx_left_in[62], chanx_left_in[103], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size6 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[20], chanx_left_in[61], chanx_left_in[102], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size6 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[19], chanx_left_in[60], chanx_left_in[101], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size6_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_11_sram_inv[0:2]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size6 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[18], chanx_left_in[59], chanx_left_in[100], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size6_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_12_sram_inv[0:2]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size6 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[17], chanx_left_in[58], chanx_left_in[99], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size6_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_13_sram_inv[0:2]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size6 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[16], chanx_left_in[57], chanx_left_in[98], chanx_left_in[139]}),
		.sram(mux_tree_tapbuf_size6_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_14_sram_inv[0:2]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size6 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[15], chanx_left_in[56], chanx_left_in[97], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size6_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_15_sram_inv[0:2]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size6 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[14], chanx_left_in[55], chanx_left_in[96], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size6_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_16_sram_inv[0:2]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size6 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[13], chanx_left_in[54], chanx_left_in[95], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size6_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_17_sram_inv[0:2]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size6 mux_top_track_232 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[12], chanx_left_in[53], chanx_left_in[94], chanx_left_in[135]}),
		.sram(mux_tree_tapbuf_size6_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_18_sram_inv[0:2]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size6 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[11], chanx_left_in[52], chanx_left_in[93], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size6_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_19_sram_inv[0:2]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size6 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[10], chanx_left_in[51], chanx_left_in[92], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size6_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_20_sram_inv[0:2]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size6 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[9], chanx_left_in[50], chanx_left_in[91], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size6_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_21_sram_inv[0:2]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size6 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[8], chanx_left_in[49], chanx_left_in[90], chanx_left_in[131]}),
		.sram(mux_tree_tapbuf_size6_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_22_sram_inv[0:2]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size6 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[7], chanx_left_in[48], chanx_left_in[89], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size6_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_23_sram_inv[0:2]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size6 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[6], chanx_left_in[47], chanx_left_in[88], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size6_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_24_sram_inv[0:2]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size6 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[5], chanx_left_in[46], chanx_left_in[87], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size6_25_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_25_sram_inv[0:2]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size6 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[4], chanx_left_in[45], chanx_left_in[86], chanx_left_in[127]}),
		.sram(mux_tree_tapbuf_size6_26_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_26_sram_inv[0:2]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size6 mux_top_track_304 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[3], chanx_left_in[44], chanx_left_in[85], chanx_left_in[126]}),
		.sram(mux_tree_tapbuf_size6_27_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_27_sram_inv[0:2]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size6 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[2], chanx_left_in[43], chanx_left_in[84], chanx_left_in[125]}),
		.sram(mux_tree_tapbuf_size6_28_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_28_sram_inv[0:2]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size6 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_left_in[1], chanx_left_in[42], chanx_left_in[83], chanx_left_in[124]}),
		.sram(mux_tree_tapbuf_size6_29_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_29_sram_inv[0:2]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size6 mux_bottom_track_1 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[1], chanx_left_in[42], chanx_left_in[83], chanx_left_in[124]}),
		.sram(mux_tree_tapbuf_size6_30_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_30_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size6 mux_bottom_track_9 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[2], chanx_left_in[43], chanx_left_in[84], chanx_left_in[125]}),
		.sram(mux_tree_tapbuf_size6_31_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_31_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size6 mux_bottom_track_17 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[3], chanx_left_in[44], chanx_left_in[85], chanx_left_in[126]}),
		.sram(mux_tree_tapbuf_size6_32_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_32_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size6 mux_bottom_track_25 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[4], chanx_left_in[45], chanx_left_in[86], chanx_left_in[127]}),
		.sram(mux_tree_tapbuf_size6_33_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_33_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size6 mux_bottom_track_33 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[5], chanx_left_in[46], chanx_left_in[87], chanx_left_in[128]}),
		.sram(mux_tree_tapbuf_size6_34_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_34_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size6 mux_bottom_track_41 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[6], chanx_left_in[47], chanx_left_in[88], chanx_left_in[129]}),
		.sram(mux_tree_tapbuf_size6_35_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_35_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size6 mux_bottom_track_49 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[7], chanx_left_in[48], chanx_left_in[89], chanx_left_in[130]}),
		.sram(mux_tree_tapbuf_size6_36_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_36_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_57 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[8], chanx_left_in[49], chanx_left_in[90], chanx_left_in[131]}),
		.sram(mux_tree_tapbuf_size6_37_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_37_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size6 mux_bottom_track_65 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[9], chanx_left_in[50], chanx_left_in[91], chanx_left_in[132]}),
		.sram(mux_tree_tapbuf_size6_38_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_38_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size6 mux_bottom_track_129 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[17], chanx_left_in[58], chanx_left_in[99], chanx_left_in[140]}),
		.sram(mux_tree_tapbuf_size6_39_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_39_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size6 mux_bottom_track_193 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[25], chanx_left_in[66], chanx_left_in[107], chanx_left_in[148]}),
		.sram(mux_tree_tapbuf_size6_40_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_40_sram_inv[0:2]),
		.out(chany_bottom_out[96]));

	mux_tree_tapbuf_size6 mux_bottom_track_257 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[33], chanx_left_in[74], chanx_left_in[115], chanx_left_in[156]}),
		.sram(mux_tree_tapbuf_size6_41_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_41_sram_inv[0:2]),
		.out(chany_bottom_out[128]));

	mux_tree_tapbuf_size6 mux_bottom_track_321 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_3_, chanx_left_in[0], chanx_left_in[41], chanx_left_in[82], chanx_left_in[123]}),
		.sram(mux_tree_tapbuf_size6_42_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_42_sram_inv[0:2]),
		.out(chany_bottom_out[160]));

	mux_tree_tapbuf_size6_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_11_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_12_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_13_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_14_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_15_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_16_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_17_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_18_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_19_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_20_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_21_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_22_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_23_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_24_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_25_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_25_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_26_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_26_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_27_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_27_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_28_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_28_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_29_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_29_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_30_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_30_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_31_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_31_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_32_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_32_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_33_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_33_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_34_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_34_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_35_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_35_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_36_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_36_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_37_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_37_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_38_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_38_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_39_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_39_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_40_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_40_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_41_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_41_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_42_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_42_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_bottom_track_73 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[10], chanx_left_in[51], chanx_left_in[92], chanx_left_in[133]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size5 mux_bottom_track_81 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[11], chanx_left_in[52], chanx_left_in[93], chanx_left_in[134]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size5 mux_bottom_track_89 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[12], chanx_left_in[53], chanx_left_in[94], chanx_left_in[135]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size5 mux_bottom_track_97 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[13], chanx_left_in[54], chanx_left_in[95], chanx_left_in[136]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size5 mux_bottom_track_105 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[14], chanx_left_in[55], chanx_left_in[96], chanx_left_in[137]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size5 mux_bottom_track_113 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[15], chanx_left_in[56], chanx_left_in[97], chanx_left_in[138]}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size5 mux_bottom_track_121 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[16], chanx_left_in[57], chanx_left_in[98], chanx_left_in[139]}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size5 mux_bottom_track_137 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[18], chanx_left_in[59], chanx_left_in[100], chanx_left_in[141]}),
		.sram(mux_tree_tapbuf_size5_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_7_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size5 mux_bottom_track_145 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[19], chanx_left_in[60], chanx_left_in[101], chanx_left_in[142]}),
		.sram(mux_tree_tapbuf_size5_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_8_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size5 mux_bottom_track_153 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[20], chanx_left_in[61], chanx_left_in[102], chanx_left_in[143]}),
		.sram(mux_tree_tapbuf_size5_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_9_sram_inv[0:2]),
		.out(chany_bottom_out[76]));

	mux_tree_tapbuf_size5 mux_bottom_track_161 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[21], chanx_left_in[62], chanx_left_in[103], chanx_left_in[144]}),
		.sram(mux_tree_tapbuf_size5_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_10_sram_inv[0:2]),
		.out(chany_bottom_out[80]));

	mux_tree_tapbuf_size5 mux_bottom_track_169 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[22], chanx_left_in[63], chanx_left_in[104], chanx_left_in[145]}),
		.sram(mux_tree_tapbuf_size5_11_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_11_sram_inv[0:2]),
		.out(chany_bottom_out[84]));

	mux_tree_tapbuf_size5 mux_bottom_track_177 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[23], chanx_left_in[64], chanx_left_in[105], chanx_left_in[146]}),
		.sram(mux_tree_tapbuf_size5_12_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_12_sram_inv[0:2]),
		.out(chany_bottom_out[88]));

	mux_tree_tapbuf_size5 mux_bottom_track_185 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[24], chanx_left_in[65], chanx_left_in[106], chanx_left_in[147]}),
		.sram(mux_tree_tapbuf_size5_13_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_13_sram_inv[0:2]),
		.out(chany_bottom_out[92]));

	mux_tree_tapbuf_size5 mux_bottom_track_201 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[26], chanx_left_in[67], chanx_left_in[108], chanx_left_in[149]}),
		.sram(mux_tree_tapbuf_size5_14_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_14_sram_inv[0:2]),
		.out(chany_bottom_out[100]));

	mux_tree_tapbuf_size5 mux_bottom_track_209 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[27], chanx_left_in[68], chanx_left_in[109], chanx_left_in[150]}),
		.sram(mux_tree_tapbuf_size5_15_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_15_sram_inv[0:2]),
		.out(chany_bottom_out[104]));

	mux_tree_tapbuf_size5 mux_bottom_track_217 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[28], chanx_left_in[69], chanx_left_in[110], chanx_left_in[151]}),
		.sram(mux_tree_tapbuf_size5_16_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_16_sram_inv[0:2]),
		.out(chany_bottom_out[108]));

	mux_tree_tapbuf_size5 mux_bottom_track_225 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[29], chanx_left_in[70], chanx_left_in[111], chanx_left_in[152]}),
		.sram(mux_tree_tapbuf_size5_17_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_17_sram_inv[0:2]),
		.out(chany_bottom_out[112]));

	mux_tree_tapbuf_size5 mux_bottom_track_233 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[30], chanx_left_in[71], chanx_left_in[112], chanx_left_in[153]}),
		.sram(mux_tree_tapbuf_size5_18_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_18_sram_inv[0:2]),
		.out(chany_bottom_out[116]));

	mux_tree_tapbuf_size5 mux_bottom_track_241 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[31], chanx_left_in[72], chanx_left_in[113], chanx_left_in[154]}),
		.sram(mux_tree_tapbuf_size5_19_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_19_sram_inv[0:2]),
		.out(chany_bottom_out[120]));

	mux_tree_tapbuf_size5 mux_bottom_track_249 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[32], chanx_left_in[73], chanx_left_in[114], chanx_left_in[155]}),
		.sram(mux_tree_tapbuf_size5_20_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_20_sram_inv[0:2]),
		.out(chany_bottom_out[124]));

	mux_tree_tapbuf_size5 mux_bottom_track_265 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_left_in[34], chanx_left_in[75], chanx_left_in[116], chanx_left_in[157]}),
		.sram(mux_tree_tapbuf_size5_21_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_21_sram_inv[0:2]),
		.out(chany_bottom_out[132]));

	mux_tree_tapbuf_size5 mux_bottom_track_273 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_left_in[35], chanx_left_in[76], chanx_left_in[117], chanx_left_in[158]}),
		.sram(mux_tree_tapbuf_size5_22_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_22_sram_inv[0:2]),
		.out(chany_bottom_out[136]));

	mux_tree_tapbuf_size5 mux_bottom_track_281 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_left_in[36], chanx_left_in[77], chanx_left_in[118], chanx_left_in[159]}),
		.sram(mux_tree_tapbuf_size5_23_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_23_sram_inv[0:2]),
		.out(chany_bottom_out[140]));

	mux_tree_tapbuf_size5 mux_bottom_track_289 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_left_in[37], chanx_left_in[78], chanx_left_in[119], chanx_left_in[160]}),
		.sram(mux_tree_tapbuf_size5_24_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_24_sram_inv[0:2]),
		.out(chany_bottom_out[144]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_7_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_9_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_10_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_11_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_11_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_12_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_12_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_13_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_13_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_14_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_14_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_15_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_15_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_16_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_16_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_17_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_17_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_18_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_18_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_19_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_19_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_20_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_20_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_21_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_21_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_22_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_22_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_23_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_23_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_24_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_24_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_bottom_track_297 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_left_in[38], chanx_left_in[79], chanx_left_in[120]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_bottom_out[148]));

	mux_tree_tapbuf_size4 mux_bottom_track_305 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_left_in[39], chanx_left_in[80], chanx_left_in[121]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_bottom_out[152]));

	mux_tree_tapbuf_size4 mux_bottom_track_313 (
		.in({bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_left_in[40], chanx_left_in[81], chanx_left_in[122]}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chany_bottom_out[156]));

	mux_tree_tapbuf_size4 mux_left_track_1 (
		.in({chany_top_in[0], chany_top_in[3], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chanx_left_out[0]));

	mux_tree_tapbuf_size4 mux_left_track_3 (
		.in({chany_bottom_in[0], chany_bottom_in[3], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_4_sram_inv[0:2]),
		.out(chanx_left_out[1]));

	mux_tree_tapbuf_size4 mux_left_track_5 (
		.in({chany_bottom_in[1], chany_bottom_in[7], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_5_sram_inv[0:2]),
		.out(chanx_left_out[2]));

	mux_tree_tapbuf_size4 mux_left_track_7 (
		.in({chany_bottom_in[2], chany_bottom_in[11], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_6_sram_inv[0:2]),
		.out(chanx_left_out[3]));

	mux_tree_tapbuf_size4 mux_left_track_9 (
		.in({chany_bottom_in[4], chany_bottom_in[15], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_7_sram_inv[0:2]),
		.out(chanx_left_out[4]));

	mux_tree_tapbuf_size4 mux_left_track_11 (
		.in({chany_bottom_in[5], chany_bottom_in[19], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_8_sram_inv[0:2]),
		.out(chanx_left_out[5]));

	mux_tree_tapbuf_size4 mux_left_track_13 (
		.in({chany_bottom_in[6], chany_bottom_in[23], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_9_sram_inv[0:2]),
		.out(chanx_left_out[6]));

	mux_tree_tapbuf_size4 mux_left_track_15 (
		.in({chany_bottom_in[8], chany_bottom_in[27], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size4_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_10_sram_inv[0:2]),
		.out(chanx_left_out[7]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_bottom_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_3 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_5 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_5_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_7 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_6_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_7_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_11 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_8_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_13 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_9_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_left_track_15 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_10_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_left_track_17 (
		.in({chany_bottom_in[9], chany_bottom_in[31], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chanx_left_out[8]));

	mux_tree_tapbuf_size3 mux_left_track_21 (
		.in({chany_bottom_in[12], chany_bottom_in[39], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chanx_left_out[10]));

	mux_tree_tapbuf_size3 mux_left_track_23 (
		.in({chany_bottom_in[13], chany_bottom_in[43], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chanx_left_out[11]));

	mux_tree_tapbuf_size3 mux_left_track_25 (
		.in({chany_bottom_in[14], chany_bottom_in[47], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chanx_left_out[12]));

	mux_tree_tapbuf_size3 mux_left_track_27 (
		.in({chany_bottom_in[16], chany_bottom_in[51], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chanx_left_out[13]));

	mux_tree_tapbuf_size3 mux_left_track_29 (
		.in({chany_bottom_in[17], chany_bottom_in[55], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chanx_left_out[14]));

	mux_tree_tapbuf_size3 mux_left_track_31 (
		.in({chany_bottom_in[18], chany_bottom_in[59], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chanx_left_out[15]));

	mux_tree_tapbuf_size3 mux_left_track_33 (
		.in({chany_bottom_in[20], chany_bottom_in[63], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chanx_left_out[16]));

	mux_tree_tapbuf_size3 mux_left_track_35 (
		.in({chany_bottom_in[21], chany_bottom_in[67], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chanx_left_out[17]));

	mux_tree_tapbuf_size3 mux_left_track_37 (
		.in({chany_bottom_in[22], chany_bottom_in[71], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chanx_left_out[18]));

	mux_tree_tapbuf_size3 mux_left_track_41 (
		.in({chany_bottom_in[25], chany_bottom_in[79], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chanx_left_out[20]));

	mux_tree_tapbuf_size3 mux_left_track_43 (
		.in({chany_bottom_in[26], chany_bottom_in[83], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chanx_left_out[21]));

	mux_tree_tapbuf_size3 mux_left_track_45 (
		.in({chany_bottom_in[28], chany_bottom_in[87], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chanx_left_out[22]));

	mux_tree_tapbuf_size3 mux_left_track_47 (
		.in({chany_bottom_in[29], chany_bottom_in[91], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chanx_left_out[23]));

	mux_tree_tapbuf_size3 mux_left_track_49 (
		.in({chany_bottom_in[30], chany_bottom_in[95], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chanx_left_out[24]));

	mux_tree_tapbuf_size3 mux_left_track_51 (
		.in({chany_bottom_in[32], chany_bottom_in[99], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chanx_left_out[25]));

	mux_tree_tapbuf_size3 mux_left_track_53 (
		.in({chany_bottom_in[33], chany_bottom_in[103], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chanx_left_out[26]));

	mux_tree_tapbuf_size3 mux_left_track_55 (
		.in({chany_bottom_in[34], chany_bottom_in[107], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chanx_left_out[27]));

	mux_tree_tapbuf_size3 mux_left_track_57 (
		.in({chany_bottom_in[36], chany_bottom_in[111], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chanx_left_out[28]));

	mux_tree_tapbuf_size3 mux_left_track_61 (
		.in({chany_bottom_in[38], chany_bottom_in[119], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chanx_left_out[30]));

	mux_tree_tapbuf_size3 mux_left_track_63 (
		.in({chany_bottom_in[40], chany_bottom_in[123], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chanx_left_out[31]));

	mux_tree_tapbuf_size3 mux_left_track_65 (
		.in({chany_bottom_in[41], chany_bottom_in[127], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chanx_left_out[32]));

	mux_tree_tapbuf_size3 mux_left_track_67 (
		.in({chany_bottom_in[42], chany_bottom_in[131], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chanx_left_out[33]));

	mux_tree_tapbuf_size3 mux_left_track_69 (
		.in({chany_bottom_in[44], chany_bottom_in[135], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chanx_left_out[34]));

	mux_tree_tapbuf_size3 mux_left_track_71 (
		.in({chany_bottom_in[45], chany_bottom_in[139], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chanx_left_out[35]));

	mux_tree_tapbuf_size3 mux_left_track_73 (
		.in({chany_bottom_in[46], chany_bottom_in[143], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chanx_left_out[36]));

	mux_tree_tapbuf_size3 mux_left_track_75 (
		.in({chany_bottom_in[48], chany_bottom_in[147], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chanx_left_out[37]));

	mux_tree_tapbuf_size3 mux_left_track_77 (
		.in({chany_bottom_in[49], chany_bottom_in[151], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chanx_left_out[38]));

	mux_tree_tapbuf_size3 mux_left_track_81 (
		.in({chany_bottom_in[52], chany_bottom_in[159], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chanx_left_out[40]));

	mux_tree_tapbuf_size3 mux_left_track_83 (
		.in({chany_bottom_in[53], chany_bottom_in[160], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chanx_left_out[41]));

	mux_tree_tapbuf_size3 mux_left_track_85 (
		.in({chany_top_in[158], chany_bottom_in[54], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chanx_left_out[42]));

	mux_tree_tapbuf_size3 mux_left_track_87 (
		.in({chany_top_in[157], chany_bottom_in[56], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chanx_left_out[43]));

	mux_tree_tapbuf_size3 mux_left_track_89 (
		.in({chany_top_in[156], chany_bottom_in[57], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chanx_left_out[44]));

	mux_tree_tapbuf_size3 mux_left_track_91 (
		.in({chany_top_in[154], chany_bottom_in[58], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chanx_left_out[45]));

	mux_tree_tapbuf_size3 mux_left_track_93 (
		.in({chany_top_in[153], chany_bottom_in[60], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chanx_left_out[46]));

	mux_tree_tapbuf_size3 mux_left_track_95 (
		.in({chany_top_in[152], chany_bottom_in[61], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chanx_left_out[47]));

	mux_tree_tapbuf_size3 mux_left_track_97 (
		.in({chany_top_in[150], chany_bottom_in[62], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chanx_left_out[48]));

	mux_tree_tapbuf_size3 mux_left_track_101 (
		.in({chany_top_in[148], chany_bottom_in[65], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chanx_left_out[50]));

	mux_tree_tapbuf_size3 mux_left_track_103 (
		.in({chany_top_in[146], chany_bottom_in[66], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chanx_left_out[51]));

	mux_tree_tapbuf_size3 mux_left_track_105 (
		.in({chany_top_in[145], chany_bottom_in[68], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chanx_left_out[52]));

	mux_tree_tapbuf_size3 mux_left_track_107 (
		.in({chany_top_in[144], chany_bottom_in[69], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chanx_left_out[53]));

	mux_tree_tapbuf_size3 mux_left_track_109 (
		.in({chany_top_in[142], chany_bottom_in[70], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chanx_left_out[54]));

	mux_tree_tapbuf_size3 mux_left_track_111 (
		.in({chany_top_in[141], chany_bottom_in[72], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chanx_left_out[55]));

	mux_tree_tapbuf_size3 mux_left_track_113 (
		.in({chany_top_in[140], chany_bottom_in[73], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chanx_left_out[56]));

	mux_tree_tapbuf_size3 mux_left_track_115 (
		.in({chany_top_in[138], chany_bottom_in[74], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chanx_left_out[57]));

	mux_tree_tapbuf_size3 mux_left_track_117 (
		.in({chany_top_in[137], chany_bottom_in[76], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chanx_left_out[58]));

	mux_tree_tapbuf_size3 mux_left_track_121 (
		.in({chany_top_in[134], chany_bottom_in[78], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chanx_left_out[60]));

	mux_tree_tapbuf_size3 mux_left_track_123 (
		.in({chany_top_in[133], chany_bottom_in[80], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chanx_left_out[61]));

	mux_tree_tapbuf_size3 mux_left_track_125 (
		.in({chany_top_in[132], chany_bottom_in[81], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chanx_left_out[62]));

	mux_tree_tapbuf_size3 mux_left_track_127 (
		.in({chany_top_in[130], chany_bottom_in[82], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chanx_left_out[63]));

	mux_tree_tapbuf_size3 mux_left_track_129 (
		.in({chany_top_in[129], chany_bottom_in[84], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chanx_left_out[64]));

	mux_tree_tapbuf_size3 mux_left_track_131 (
		.in({chany_top_in[128], chany_bottom_in[85], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chanx_left_out[65]));

	mux_tree_tapbuf_size3 mux_left_track_133 (
		.in({chany_top_in[126], chany_bottom_in[86], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chanx_left_out[66]));

	mux_tree_tapbuf_size3 mux_left_track_135 (
		.in({chany_top_in[125], chany_bottom_in[88], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chanx_left_out[67]));

	mux_tree_tapbuf_size3 mux_left_track_137 (
		.in({chany_top_in[124], chany_bottom_in[89], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chanx_left_out[68]));

	mux_tree_tapbuf_size3 mux_left_track_141 (
		.in({chany_top_in[121], chany_bottom_in[92], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chanx_left_out[70]));

	mux_tree_tapbuf_size3 mux_left_track_143 (
		.in({chany_top_in[120], chany_bottom_in[93], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chanx_left_out[71]));

	mux_tree_tapbuf_size3 mux_left_track_145 (
		.in({chany_top_in[118], chany_bottom_in[94], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chanx_left_out[72]));

	mux_tree_tapbuf_size3 mux_left_track_147 (
		.in({chany_top_in[117], chany_bottom_in[96], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chanx_left_out[73]));

	mux_tree_tapbuf_size3 mux_left_track_149 (
		.in({chany_top_in[116], chany_bottom_in[97], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chanx_left_out[74]));

	mux_tree_tapbuf_size3 mux_left_track_151 (
		.in({chany_top_in[114], chany_bottom_in[98], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_60_sram_inv[0:1]),
		.out(chanx_left_out[75]));

	mux_tree_tapbuf_size3 mux_left_track_153 (
		.in({chany_top_in[113], chany_bottom_in[100], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_61_sram_inv[0:1]),
		.out(chanx_left_out[76]));

	mux_tree_tapbuf_size3 mux_left_track_155 (
		.in({chany_top_in[112], chany_bottom_in[101], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_62_sram_inv[0:1]),
		.out(chanx_left_out[77]));

	mux_tree_tapbuf_size3 mux_left_track_157 (
		.in({chany_top_in[110], chany_bottom_in[102], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_63_sram_inv[0:1]),
		.out(chanx_left_out[78]));

	mux_tree_tapbuf_size3 mux_left_track_161 (
		.in({chany_top_in[108], chany_bottom_in[105], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_64_sram_inv[0:1]),
		.out(chanx_left_out[80]));

	mux_tree_tapbuf_size3 mux_left_track_163 (
		.in({chany_top_in[106], chany_bottom_in[106], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_65_sram_inv[0:1]),
		.out(chanx_left_out[81]));

	mux_tree_tapbuf_size3 mux_left_track_165 (
		.in({chany_top_in[105], chany_bottom_in[108], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_66_sram_inv[0:1]),
		.out(chanx_left_out[82]));

	mux_tree_tapbuf_size3 mux_left_track_167 (
		.in({chany_top_in[104], chany_bottom_in[109], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_67_sram_inv[0:1]),
		.out(chanx_left_out[83]));

	mux_tree_tapbuf_size3 mux_left_track_169 (
		.in({chany_top_in[102], chany_bottom_in[110], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_68_sram_inv[0:1]),
		.out(chanx_left_out[84]));

	mux_tree_tapbuf_size3 mux_left_track_171 (
		.in({chany_top_in[101], chany_bottom_in[112], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_69_sram_inv[0:1]),
		.out(chanx_left_out[85]));

	mux_tree_tapbuf_size3 mux_left_track_173 (
		.in({chany_top_in[100], chany_bottom_in[113], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_70_sram_inv[0:1]),
		.out(chanx_left_out[86]));

	mux_tree_tapbuf_size3 mux_left_track_175 (
		.in({chany_top_in[98], chany_bottom_in[114], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_71_sram_inv[0:1]),
		.out(chanx_left_out[87]));

	mux_tree_tapbuf_size3 mux_left_track_177 (
		.in({chany_top_in[97], chany_bottom_in[116], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_72_sram_inv[0:1]),
		.out(chanx_left_out[88]));

	mux_tree_tapbuf_size3 mux_left_track_181 (
		.in({chany_top_in[94], chany_bottom_in[118], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_73_sram_inv[0:1]),
		.out(chanx_left_out[90]));

	mux_tree_tapbuf_size3 mux_left_track_183 (
		.in({chany_top_in[93], chany_bottom_in[120], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_74_sram_inv[0:1]),
		.out(chanx_left_out[91]));

	mux_tree_tapbuf_size3 mux_left_track_185 (
		.in({chany_top_in[92], chany_bottom_in[121], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_75_sram_inv[0:1]),
		.out(chanx_left_out[92]));

	mux_tree_tapbuf_size3 mux_left_track_187 (
		.in({chany_top_in[90], chany_bottom_in[122], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_76_sram_inv[0:1]),
		.out(chanx_left_out[93]));

	mux_tree_tapbuf_size3 mux_left_track_189 (
		.in({chany_top_in[89], chany_bottom_in[124], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_77_sram_inv[0:1]),
		.out(chanx_left_out[94]));

	mux_tree_tapbuf_size3 mux_left_track_191 (
		.in({chany_top_in[88], chany_bottom_in[125], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_78_sram_inv[0:1]),
		.out(chanx_left_out[95]));

	mux_tree_tapbuf_size3 mux_left_track_193 (
		.in({chany_top_in[86], chany_bottom_in[126], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_79_sram_inv[0:1]),
		.out(chanx_left_out[96]));

	mux_tree_tapbuf_size3 mux_left_track_195 (
		.in({chany_top_in[85], chany_bottom_in[128], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_80_sram_inv[0:1]),
		.out(chanx_left_out[97]));

	mux_tree_tapbuf_size3 mux_left_track_197 (
		.in({chany_top_in[84], chany_bottom_in[129], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_81_sram_inv[0:1]),
		.out(chanx_left_out[98]));

	mux_tree_tapbuf_size3 mux_left_track_201 (
		.in({chany_top_in[81], chany_bottom_in[132], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_82_sram_inv[0:1]),
		.out(chanx_left_out[100]));

	mux_tree_tapbuf_size3 mux_left_track_203 (
		.in({chany_top_in[80], chany_bottom_in[133], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_83_sram_inv[0:1]),
		.out(chanx_left_out[101]));

	mux_tree_tapbuf_size3 mux_left_track_205 (
		.in({chany_top_in[78], chany_bottom_in[134], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_84_sram_inv[0:1]),
		.out(chanx_left_out[102]));

	mux_tree_tapbuf_size3 mux_left_track_207 (
		.in({chany_top_in[77], chany_bottom_in[136], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_85_sram_inv[0:1]),
		.out(chanx_left_out[103]));

	mux_tree_tapbuf_size3 mux_left_track_209 (
		.in({chany_top_in[76], chany_bottom_in[137], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_86_sram_inv[0:1]),
		.out(chanx_left_out[104]));

	mux_tree_tapbuf_size3 mux_left_track_211 (
		.in({chany_top_in[74], chany_bottom_in[138], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_87_sram_inv[0:1]),
		.out(chanx_left_out[105]));

	mux_tree_tapbuf_size3 mux_left_track_213 (
		.in({chany_top_in[73], chany_bottom_in[140], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_88_sram_inv[0:1]),
		.out(chanx_left_out[106]));

	mux_tree_tapbuf_size3 mux_left_track_215 (
		.in({chany_top_in[72], chany_bottom_in[141], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_89_sram_inv[0:1]),
		.out(chanx_left_out[107]));

	mux_tree_tapbuf_size3 mux_left_track_217 (
		.in({chany_top_in[70], chany_bottom_in[142], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_90_sram_inv[0:1]),
		.out(chanx_left_out[108]));

	mux_tree_tapbuf_size3 mux_left_track_221 (
		.in({chany_top_in[68], chany_bottom_in[145], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_91_sram_inv[0:1]),
		.out(chanx_left_out[110]));

	mux_tree_tapbuf_size3 mux_left_track_223 (
		.in({chany_top_in[66], chany_bottom_in[146], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_92_sram_inv[0:1]),
		.out(chanx_left_out[111]));

	mux_tree_tapbuf_size3 mux_left_track_225 (
		.in({chany_top_in[65], chany_bottom_in[148], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_93_sram_inv[0:1]),
		.out(chanx_left_out[112]));

	mux_tree_tapbuf_size3 mux_left_track_227 (
		.in({chany_top_in[64], chany_bottom_in[149], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_94_sram_inv[0:1]),
		.out(chanx_left_out[113]));

	mux_tree_tapbuf_size3 mux_left_track_229 (
		.in({chany_top_in[62], chany_bottom_in[150], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_95_sram_inv[0:1]),
		.out(chanx_left_out[114]));

	mux_tree_tapbuf_size3 mux_left_track_231 (
		.in({chany_top_in[61], chany_bottom_in[152], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_96_sram_inv[0:1]),
		.out(chanx_left_out[115]));

	mux_tree_tapbuf_size3 mux_left_track_233 (
		.in({chany_top_in[60], chany_bottom_in[153], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_97_sram_inv[0:1]),
		.out(chanx_left_out[116]));

	mux_tree_tapbuf_size3 mux_left_track_235 (
		.in({chany_top_in[58], chany_bottom_in[154], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_98_sram_inv[0:1]),
		.out(chanx_left_out[117]));

	mux_tree_tapbuf_size3 mux_left_track_237 (
		.in({chany_top_in[57], chany_bottom_in[156], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_99_sram_inv[0:1]),
		.out(chanx_left_out[118]));

	mux_tree_tapbuf_size3 mux_left_track_241 (
		.in({chany_top_in[54], chany_bottom_in[158], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_100_sram_inv[0:1]),
		.out(chanx_left_out[120]));

	mux_tree_tapbuf_size3 mux_left_track_243 (
		.in({chany_top_in[53], chany_top_in[160], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_101_sram_inv[0:1]),
		.out(chanx_left_out[121]));

	mux_tree_tapbuf_size3 mux_left_track_245 (
		.in({chany_top_in[52], chany_top_in[159], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_102_sram_inv[0:1]),
		.out(chanx_left_out[122]));

	mux_tree_tapbuf_size3 mux_left_track_247 (
		.in({chany_top_in[50], chany_top_in[155], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_103_sram_inv[0:1]),
		.out(chanx_left_out[123]));

	mux_tree_tapbuf_size3 mux_left_track_249 (
		.in({chany_top_in[49], chany_top_in[151], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_104_sram_inv[0:1]),
		.out(chanx_left_out[124]));

	mux_tree_tapbuf_size3 mux_left_track_251 (
		.in({chany_top_in[48], chany_top_in[147], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_105_sram_inv[0:1]),
		.out(chanx_left_out[125]));

	mux_tree_tapbuf_size3 mux_left_track_253 (
		.in({chany_top_in[46], chany_top_in[143], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_106_sram_inv[0:1]),
		.out(chanx_left_out[126]));

	mux_tree_tapbuf_size3 mux_left_track_255 (
		.in({chany_top_in[45], chany_top_in[139], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_107_sram_inv[0:1]),
		.out(chanx_left_out[127]));

	mux_tree_tapbuf_size3 mux_left_track_257 (
		.in({chany_top_in[44], chany_top_in[135], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_108_sram_inv[0:1]),
		.out(chanx_left_out[128]));

	mux_tree_tapbuf_size3 mux_left_track_261 (
		.in({chany_top_in[41], chany_top_in[127], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_109_sram_inv[0:1]),
		.out(chanx_left_out[130]));

	mux_tree_tapbuf_size3 mux_left_track_263 (
		.in({chany_top_in[40], chany_top_in[123], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_110_sram_inv[0:1]),
		.out(chanx_left_out[131]));

	mux_tree_tapbuf_size3 mux_left_track_265 (
		.in({chany_top_in[38], chany_top_in[119], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_111_sram_inv[0:1]),
		.out(chanx_left_out[132]));

	mux_tree_tapbuf_size3 mux_left_track_267 (
		.in({chany_top_in[37], chany_top_in[115], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_112_sram_inv[0:1]),
		.out(chanx_left_out[133]));

	mux_tree_tapbuf_size3 mux_left_track_269 (
		.in({chany_top_in[36], chany_top_in[111], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_113_sram_inv[0:1]),
		.out(chanx_left_out[134]));

	mux_tree_tapbuf_size3 mux_left_track_271 (
		.in({chany_top_in[34], chany_top_in[107], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_114_sram_inv[0:1]),
		.out(chanx_left_out[135]));

	mux_tree_tapbuf_size3 mux_left_track_273 (
		.in({chany_top_in[33], chany_top_in[103], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_115_sram_inv[0:1]),
		.out(chanx_left_out[136]));

	mux_tree_tapbuf_size3 mux_left_track_275 (
		.in({chany_top_in[32], chany_top_in[99], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_116_sram_inv[0:1]),
		.out(chanx_left_out[137]));

	mux_tree_tapbuf_size3 mux_left_track_277 (
		.in({chany_top_in[30], chany_top_in[95], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_117_sram_inv[0:1]),
		.out(chanx_left_out[138]));

	mux_tree_tapbuf_size3 mux_left_track_281 (
		.in({chany_top_in[28], chany_top_in[87], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_118_sram_inv[0:1]),
		.out(chanx_left_out[140]));

	mux_tree_tapbuf_size3 mux_left_track_283 (
		.in({chany_top_in[26], chany_top_in[83], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_119_sram_inv[0:1]),
		.out(chanx_left_out[141]));

	mux_tree_tapbuf_size3 mux_left_track_285 (
		.in({chany_top_in[25], chany_top_in[79], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_120_sram_inv[0:1]),
		.out(chanx_left_out[142]));

	mux_tree_tapbuf_size3 mux_left_track_287 (
		.in({chany_top_in[24], chany_top_in[75], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_121_sram_inv[0:1]),
		.out(chanx_left_out[143]));

	mux_tree_tapbuf_size3 mux_left_track_289 (
		.in({chany_top_in[22], chany_top_in[71], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_122_sram_inv[0:1]),
		.out(chanx_left_out[144]));

	mux_tree_tapbuf_size3 mux_left_track_291 (
		.in({chany_top_in[21], chany_top_in[67], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_123_sram_inv[0:1]),
		.out(chanx_left_out[145]));

	mux_tree_tapbuf_size3 mux_left_track_293 (
		.in({chany_top_in[20], chany_top_in[63], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_124_sram_inv[0:1]),
		.out(chanx_left_out[146]));

	mux_tree_tapbuf_size3 mux_left_track_295 (
		.in({chany_top_in[18], chany_top_in[59], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_125_sram_inv[0:1]),
		.out(chanx_left_out[147]));

	mux_tree_tapbuf_size3 mux_left_track_297 (
		.in({chany_top_in[17], chany_top_in[55], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_126_sram_inv[0:1]),
		.out(chanx_left_out[148]));

	mux_tree_tapbuf_size3 mux_left_track_301 (
		.in({chany_top_in[14], chany_top_in[47], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_127_sram_inv[0:1]),
		.out(chanx_left_out[150]));

	mux_tree_tapbuf_size3 mux_left_track_303 (
		.in({chany_top_in[13], chany_top_in[43], left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_128_sram_inv[0:1]),
		.out(chanx_left_out[151]));

	mux_tree_tapbuf_size3 mux_left_track_305 (
		.in({chany_top_in[12], chany_top_in[39], left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_129_sram_inv[0:1]),
		.out(chanx_left_out[152]));

	mux_tree_tapbuf_size3 mux_left_track_307 (
		.in({chany_top_in[10], chany_top_in[35], left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_130_sram_inv[0:1]),
		.out(chanx_left_out[153]));

	mux_tree_tapbuf_size3 mux_left_track_309 (
		.in({chany_top_in[9], chany_top_in[31], left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_131_sram_inv[0:1]),
		.out(chanx_left_out[154]));

	mux_tree_tapbuf_size3 mux_left_track_311 (
		.in({chany_top_in[8], chany_top_in[27], left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_132_sram_inv[0:1]),
		.out(chanx_left_out[155]));

	mux_tree_tapbuf_size3 mux_left_track_313 (
		.in({chany_top_in[6], chany_top_in[23], left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_133_sram_inv[0:1]),
		.out(chanx_left_out[156]));

	mux_tree_tapbuf_size3 mux_left_track_315 (
		.in({chany_top_in[5], chany_top_in[19], left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_134_sram_inv[0:1]),
		.out(chanx_left_out[157]));

	mux_tree_tapbuf_size3 mux_left_track_317 (
		.in({chany_top_in[4], chany_top_in[15], left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_135_sram_inv[0:1]),
		.out(chanx_left_out[158]));

	mux_tree_tapbuf_size3 mux_left_track_321 (
		.in({chany_top_in[1], chany_top_in[7], left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_136_sram_inv[0:1]),
		.out(chanx_left_out[160]));

	mux_tree_tapbuf_size3_mem mem_left_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_21 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_23 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_27 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_29 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_31 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_35 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_37 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_43 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_45 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_47 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_51 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_53 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_55 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_61 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_63 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_67 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_69 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_71 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_75 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_77 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_83 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_85 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_87 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_91 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_93 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_95 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_101 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_103 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_107 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_109 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_111 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_115 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_117 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_123 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_125 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_127 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_131 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_133 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_135 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_141 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_143 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_147 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_149 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_151 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_60_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_153 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_61_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_155 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_62_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_157 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_63_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_161 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_64_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_163 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_65_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_165 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_66_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_167 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_67_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_169 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_68_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_171 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_69_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_173 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_70_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_175 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_71_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_177 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_72_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_181 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_73_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_183 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_74_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_185 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_75_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_187 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_76_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_189 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_77_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_191 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_78_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_193 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_79_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_195 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_80_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_197 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_81_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_201 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_82_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_203 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_83_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_205 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_84_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_207 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_85_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_209 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_86_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_211 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_87_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_213 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_88_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_215 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_89_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_217 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_90_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_221 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_91_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_223 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_92_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_225 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_93_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_227 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_94_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_229 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_95_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_231 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_96_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_233 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_97_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_235 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_98_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_237 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_99_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_241 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_100_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_243 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_101_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_245 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_102_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_247 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_103_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_249 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_104_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_251 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_105_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_253 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_106_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_255 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_107_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_257 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_108_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_261 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_109_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_263 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_110_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_265 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_111_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_267 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_112_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_269 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_113_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_271 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_114_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_273 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_115_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_275 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_116_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_277 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_117_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_281 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_118_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_283 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_119_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_285 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_120_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_287 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_121_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_289 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_122_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_291 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_123_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_293 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_124_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_295 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_125_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_297 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_126_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_301 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_127_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_303 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_128_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_305 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_129_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_307 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_130_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_309 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_131_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_311 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_132_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_313 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_133_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_315 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_134_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_317 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_135_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_left_track_321 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_136_sram_inv[0:1]));

	mux_tree_tapbuf_size2 mux_left_track_19 (
		.in({chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chanx_left_out[9]));

	mux_tree_tapbuf_size2 mux_left_track_39 (
		.in({chany_bottom_in[24], chany_bottom_in[75]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chanx_left_out[19]));

	mux_tree_tapbuf_size2 mux_left_track_59 (
		.in({chany_bottom_in[37], chany_bottom_in[115]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chanx_left_out[29]));

	mux_tree_tapbuf_size2 mux_left_track_79 (
		.in({chany_bottom_in[50], chany_bottom_in[155]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chanx_left_out[39]));

	mux_tree_tapbuf_size2 mux_left_track_99 (
		.in({chany_top_in[149], chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chanx_left_out[49]));

	mux_tree_tapbuf_size2 mux_left_track_119 (
		.in({chany_top_in[136], chany_bottom_in[77]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chanx_left_out[59]));

	mux_tree_tapbuf_size2 mux_left_track_139 (
		.in({chany_top_in[122], chany_bottom_in[90]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chanx_left_out[69]));

	mux_tree_tapbuf_size2 mux_left_track_159 (
		.in({chany_top_in[109], chany_bottom_in[104]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chanx_left_out[79]));

	mux_tree_tapbuf_size2 mux_left_track_179 (
		.in({chany_top_in[96], chany_bottom_in[117]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chanx_left_out[89]));

	mux_tree_tapbuf_size2 mux_left_track_199 (
		.in({chany_top_in[82], chany_bottom_in[130]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chanx_left_out[99]));

	mux_tree_tapbuf_size2 mux_left_track_219 (
		.in({chany_top_in[69], chany_bottom_in[144]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chanx_left_out[109]));

	mux_tree_tapbuf_size2 mux_left_track_239 (
		.in({chany_top_in[56], chany_bottom_in[157]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chanx_left_out[119]));

	mux_tree_tapbuf_size2 mux_left_track_259 (
		.in({chany_top_in[42], chany_top_in[131]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chanx_left_out[129]));

	mux_tree_tapbuf_size2 mux_left_track_279 (
		.in({chany_top_in[29], chany_top_in[91]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chanx_left_out[139]));

	mux_tree_tapbuf_size2 mux_left_track_299 (
		.in({chany_top_in[16], chany_top_in[51]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chanx_left_out[149]));

	mux_tree_tapbuf_size2 mux_left_track_319 (
		.in({chany_top_in[2], chany_top_in[11]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chanx_left_out[159]));

	mux_tree_tapbuf_size2_mem mem_left_track_19 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_39 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_59 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_79 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_99 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_119 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_139 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_159 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_179 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_199 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_219 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_239 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_259 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_279 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_299 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_left_track_319 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_18__16_ -----

//----- Default net type -----
`default_nettype wire



