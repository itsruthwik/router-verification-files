//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][2]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Jun 29 10:24:45 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__2_ -----
module sb_0__2_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:72] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:72] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_;
//----- INPUT PORTS -----
input [0:72] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:72] chany_top_out;
//----- OUTPUT PORTS -----
output [0:72] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:72] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_1_sram;
wire [0:3] mux_tree_tapbuf_size10_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size10_2_sram;
wire [0:3] mux_tree_tapbuf_size10_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size10_mem_2_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_11_sram;
wire [0:3] mux_tree_tapbuf_size11_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_12_sram;
wire [0:3] mux_tree_tapbuf_size11_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_13_sram;
wire [0:3] mux_tree_tapbuf_size11_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_10_sram;
wire [0:3] mux_tree_tapbuf_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_11_sram;
wire [0:3] mux_tree_tapbuf_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_12_sram;
wire [0:3] mux_tree_tapbuf_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_13_sram;
wire [0:3] mux_tree_tapbuf_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_14_sram;
wire [0:3] mux_tree_tapbuf_size13_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_15_sram;
wire [0:3] mux_tree_tapbuf_size13_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_16_sram;
wire [0:3] mux_tree_tapbuf_size13_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_17_sram;
wire [0:3] mux_tree_tapbuf_size13_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_18_sram;
wire [0:3] mux_tree_tapbuf_size13_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_9_sram;
wire [0:3] mux_tree_tapbuf_size13_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:4] mux_tree_tapbuf_size20_0_sram;
wire [0:4] mux_tree_tapbuf_size20_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_1_sram;
wire [0:4] mux_tree_tapbuf_size20_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_2_sram;
wire [0:4] mux_tree_tapbuf_size20_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_3_sram;
wire [0:4] mux_tree_tapbuf_size20_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_4_sram;
wire [0:4] mux_tree_tapbuf_size20_4_sram_inv;
wire [0:0] mux_tree_tapbuf_size20_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_4_ccff_tail;
wire [0:4] mux_tree_tapbuf_size21_0_sram;
wire [0:4] mux_tree_tapbuf_size21_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_10_sram;
wire [0:4] mux_tree_tapbuf_size21_10_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_11_sram;
wire [0:4] mux_tree_tapbuf_size21_11_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_1_sram;
wire [0:4] mux_tree_tapbuf_size21_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_2_sram;
wire [0:4] mux_tree_tapbuf_size21_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_3_sram;
wire [0:4] mux_tree_tapbuf_size21_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_4_sram;
wire [0:4] mux_tree_tapbuf_size21_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_5_sram;
wire [0:4] mux_tree_tapbuf_size21_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_6_sram;
wire [0:4] mux_tree_tapbuf_size21_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_7_sram;
wire [0:4] mux_tree_tapbuf_size21_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_8_sram;
wire [0:4] mux_tree_tapbuf_size21_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_9_sram;
wire [0:4] mux_tree_tapbuf_size21_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size21_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size22_0_sram;
wire [0:4] mux_tree_tapbuf_size22_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_1_sram;
wire [0:4] mux_tree_tapbuf_size22_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size22_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_1_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_1_sram;
wire [0:2] mux_tree_tapbuf_size7_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size7_2_sram;
wire [0:2] mux_tree_tapbuf_size7_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size7_mem_2_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 243 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 244 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 245 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 247 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 248 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 249 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 251 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 252 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 253 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 255 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 256 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 257 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 259 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 260 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 261 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 263 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 264 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 265 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 267 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 268 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 269 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 271 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 272 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 273 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 275 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 276 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 277 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 279 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 280 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 281 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 283 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 284 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 285 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 287 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 288 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 289 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 291 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 292 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 293 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 295 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 296 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 297 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 299 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 300 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 301 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 303 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 304 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 305 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 307 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 308 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 309 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 311 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 312 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 313 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size7 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[1], chanx_right_in[20], chanx_right_in[39], chanx_right_in[58]}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size7 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[7], chanx_right_in[26], chanx_right_in[45], chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_size7_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_1_sram_inv[0:2]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size7 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[46], chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_size7_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_2_sram_inv[0:2]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size7_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_1_sram_inv[0:2]));

	mux_tree_tapbuf_size7_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[2], chanx_right_in[21], chanx_right_in[40], chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size6 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[3], chanx_right_in[22], chanx_right_in[41], chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size6 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[4], chanx_right_in[23], chanx_right_in[42], chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size6 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[5], chanx_right_in[24], chanx_right_in[43], chanx_right_in[62]}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size6 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[6], chanx_right_in[25], chanx_right_in[44], chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size6 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[9], chanx_right_in[28], chanx_right_in[47], chanx_right_in[66]}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size6 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[13], chanx_right_in[32], chanx_right_in[51], chanx_right_in[70]}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size6 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[14], chanx_right_in[33], chanx_right_in[52], chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size6 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[0], chanx_right_in[19], chanx_right_in[38], chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size6_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[10], chanx_right_in[29], chanx_right_in[48], chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size5 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[11], chanx_right_in[30], chanx_right_in[49], chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size5 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[12], chanx_right_in[31], chanx_right_in[50], chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size5 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[15], chanx_right_in[34], chanx_right_in[53], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size5 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, chanx_right_in[18], chanx_right_in[37], chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size5_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size4 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[16], chanx_right_in[35], chanx_right_in[54]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size4 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[17], chanx_right_in[36], chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size4_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size10 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size10 mux_right_track_70 (
		.in({chany_top_in[45], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_size10_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_1_sram_inv[0:3]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size10 mux_right_track_144 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size10_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_2_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size10_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_1_sram_inv[0:3]));

	mux_tree_tapbuf_size10_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size13 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size13 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size13 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size13 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size13 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size13 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size13 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size13 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size13 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, chany_bottom_in[70]}),
		.sram(mux_tree_tapbuf_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_9_sram_inv[0:3]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size13 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[72], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_10_sram_inv[0:3]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size13 mux_right_track_44 (
		.in({chany_top_in[28], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_11_sram_inv[0:3]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size13 mux_right_track_48 (
		.in({chany_top_in[30], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_12_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size13 mux_right_track_62 (
		.in({chany_top_in[40], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_13_sram_inv[0:3]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size13 mux_right_track_80 (
		.in({chany_top_in[52], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_size13_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_14_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size13 mux_right_track_98 (
		.in({chany_top_in[64], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[29]}),
		.sram(mux_tree_tapbuf_size13_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_15_sram_inv[0:3]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size13 mux_right_track_108 (
		.in({chany_top_in[70], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_size13_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_16_sram_inv[0:3]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size13 mux_right_track_116 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size13_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_17_sram_inv[0:3]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size13 mux_right_track_134 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_, chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size13_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_18_sram_inv[0:3]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size13_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_14_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_15_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_16_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_17_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size12 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size12 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size12 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size12 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size12 mux_right_track_40 (
		.in({chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size12 mux_right_track_42 (
		.in({chany_top_in[26], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, chany_bottom_in[66]}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size12 mux_right_track_46 (
		.in({chany_top_in[29], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size12 mux_right_track_54 (
		.in({chany_top_in[34], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, chany_bottom_in[58]}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size12 mux_right_track_56 (
		.in({chany_top_in[36], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size12 mux_right_track_58 (
		.in({chany_top_in[37], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size12 mux_right_track_60 (
		.in({chany_top_in[38], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size12 mux_right_track_64 (
		.in({chany_top_in[41], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size12 mux_right_track_68 (
		.in({chany_top_in[44], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size12 mux_right_track_72 (
		.in({chany_top_in[46], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, chany_bottom_in[46]}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size12 mux_right_track_74 (
		.in({chany_top_in[48], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size12 mux_right_track_76 (
		.in({chany_top_in[49], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size12 mux_right_track_78 (
		.in({chany_top_in[50], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size12 mux_right_track_82 (
		.in({chany_top_in[53], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, chany_bottom_in[40]}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size12 mux_right_track_84 (
		.in({chany_top_in[54], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size12 mux_right_track_92 (
		.in({chany_top_in[60], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size12 mux_right_track_94 (
		.in({chany_top_in[61], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size12 mux_right_track_96 (
		.in({chany_top_in[62], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, chany_bottom_in[30]}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size12 mux_right_track_100 (
		.in({chany_top_in[65], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, chany_bottom_in[28]}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size12 mux_right_track_102 (
		.in({chany_top_in[66], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, chany_bottom_in[26]}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size12 mux_right_track_104 (
		.in({chany_top_in[68], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, chany_bottom_in[25]}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size12 mux_right_track_112 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size12 mux_right_track_114 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_106_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_146_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_, chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size12 mux_right_track_118 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size12 mux_right_track_120 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size12 mux_right_track_122 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size12 mux_right_track_128 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_214_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_254_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size12 mux_right_track_132 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_46_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_82_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size12 mux_right_track_136 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_18_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_54_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_90_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_322_, chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size12 mux_right_track_138 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_286_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_326_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size12 mux_right_track_140 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_290_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_330_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size12_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size14 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_10_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_14_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_50_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_86_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_2_}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size14_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size11 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_118_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_158_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_198_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_238_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_278_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_318_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size11 mux_right_track_50 (
		.in({chany_top_in[32], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_110_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_150_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size11 mux_right_track_52 (
		.in({chany_top_in[33], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_102_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_114_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_154_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_194_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_234_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_274_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_314_, chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size11 mux_right_track_66 (
		.in({chany_top_in[42], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_22_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_58_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_94_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_142_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size11 mux_right_track_86 (
		.in({chany_top_in[56], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_26_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_62_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_98_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_182_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size11 mux_right_track_88 (
		.in({chany_top_in[57], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_134_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_174_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_186_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_226_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_266_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_306_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_6_, chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size11 mux_right_track_90 (
		.in({chany_top_in[58], right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_190_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size11 mux_right_track_106 (
		.in({chany_top_in[69], right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_222_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, chany_bottom_in[24], chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size11 mux_right_track_110 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_2_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_38_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_74_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_230_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size11 mux_right_track_124 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_126_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_166_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_206_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_246_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_298_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_338_, chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size11 mux_right_track_126 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_34_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_70_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_130_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_170_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_210_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_250_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_262_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_302_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size11_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_11_sram_inv[0:3]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size11 mux_right_track_130 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_6_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_42_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_78_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_138_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_178_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_218_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_258_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_270_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_310_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size11_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_12_sram_inv[0:3]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size11 mux_right_track_142 (
		.in({right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_30_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_66_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_122_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_162_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_202_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_242_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_282_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_294_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_channel_out_op_334_, chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_size11_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_13_sram_inv[0:3]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size11_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_11_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_12_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_13_sram_inv[0:3]));

	mux_tree_tapbuf_size21 mux_bottom_track_1 (
		.in({chanx_right_in[17], chanx_right_in[36], chanx_right_in[55], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_0_sram_inv[0:4]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size21 mux_bottom_track_17 (
		.in({chanx_right_in[15], chanx_right_in[34], chanx_right_in[53], chanx_right_in[72], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_1_sram_inv[0:4]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size21 mux_bottom_track_41 (
		.in({chanx_right_in[12], chanx_right_in[31], chanx_right_in[50], chanx_right_in[69], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_2_sram_inv[0:4]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size21 mux_bottom_track_57 (
		.in({chanx_right_in[10], chanx_right_in[29], chanx_right_in[48], chanx_right_in[67], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_3_sram_inv[0:4]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size21 mux_bottom_track_65 (
		.in({chanx_right_in[9], chanx_right_in[28], chanx_right_in[47], chanx_right_in[66], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_4_sram_inv[0:4]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size21 mux_bottom_track_73 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[46], chanx_right_in[65], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_5_sram_inv[0:4]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size21 mux_bottom_track_81 (
		.in({chanx_right_in[7], chanx_right_in[26], chanx_right_in[45], chanx_right_in[64], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_6_sram_inv[0:4]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size21 mux_bottom_track_89 (
		.in({chanx_right_in[6], chanx_right_in[25], chanx_right_in[44], chanx_right_in[63], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_7_sram_inv[0:4]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size21 mux_bottom_track_121 (
		.in({chanx_right_in[2], chanx_right_in[21], chanx_right_in[40], chanx_right_in[59], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_8_sram_inv[0:4]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size21 mux_bottom_track_129 (
		.in({chanx_right_in[1], chanx_right_in[20], chanx_right_in[39], chanx_right_in[58], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_9_sram_inv[0:4]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size21 mux_bottom_track_137 (
		.in({chanx_right_in[0], chanx_right_in[19], chanx_right_in[38], chanx_right_in[57], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_10_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_10_sram_inv[0:4]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size21 mux_bottom_track_145 (
		.in({chanx_right_in[18], chanx_right_in[37], chanx_right_in[56], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size21_11_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_11_sram_inv[0:4]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_0_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_1_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_2_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_3_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_4_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_5_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_6_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_7_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_8_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_9_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_10_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_10_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_10_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_11_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_11_sram_inv[0:4]));

	mux_tree_tapbuf_size20 mux_bottom_track_9 (
		.in({chanx_right_in[16], chanx_right_in[35], chanx_right_in[54], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size20_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_0_sram_inv[0:4]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size20 mux_bottom_track_25 (
		.in({chanx_right_in[14], chanx_right_in[33], chanx_right_in[52], chanx_right_in[71], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size20_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_1_sram_inv[0:4]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size20 mux_bottom_track_33 (
		.in({chanx_right_in[13], chanx_right_in[32], chanx_right_in[51], chanx_right_in[70], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size20_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_2_sram_inv[0:4]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size20 mux_bottom_track_105 (
		.in({chanx_right_in[4], chanx_right_in[23], chanx_right_in[42], chanx_right_in[61], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size20_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_3_sram_inv[0:4]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size20 mux_bottom_track_113 (
		.in({chanx_right_in[3], chanx_right_in[22], chanx_right_in[41], chanx_right_in[60], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size20_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_4_sram_inv[0:4]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_0_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_1_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_2_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_3_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_4_sram_inv[0:4]));

	mux_tree_tapbuf_size22 mux_bottom_track_49 (
		.in({chanx_right_in[11], chanx_right_in[30], chanx_right_in[49], chanx_right_in[68], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size22_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_0_sram_inv[0:4]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size22 mux_bottom_track_97 (
		.in({chanx_right_in[5], chanx_right_in[24], chanx_right_in[43], chanx_right_in[62], bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, bottom_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size22_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_1_sram_inv[0:4]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_0_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_1_sram_inv[0:4]));

endmodule
// ----- END Verilog module for sb_0__2_ -----

//----- Default net type -----
`default_nettype wire



