//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][0]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Fri Jul  5 01:26:08 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__0_ -----
module sb_0__0_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_,
                right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_,
                right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:284] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:284] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:284] chany_top_out;
//----- OUTPUT PORTS -----
output [0:284] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:1] mux_tree_tapbuf_size2_0_sram;
wire [0:1] mux_tree_tapbuf_size2_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_100_sram;
wire [0:1] mux_tree_tapbuf_size2_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_101_sram;
wire [0:1] mux_tree_tapbuf_size2_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_102_sram;
wire [0:1] mux_tree_tapbuf_size2_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_103_sram;
wire [0:1] mux_tree_tapbuf_size2_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_104_sram;
wire [0:1] mux_tree_tapbuf_size2_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_105_sram;
wire [0:1] mux_tree_tapbuf_size2_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_106_sram;
wire [0:1] mux_tree_tapbuf_size2_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_107_sram;
wire [0:1] mux_tree_tapbuf_size2_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_108_sram;
wire [0:1] mux_tree_tapbuf_size2_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_109_sram;
wire [0:1] mux_tree_tapbuf_size2_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_10_sram;
wire [0:1] mux_tree_tapbuf_size2_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_110_sram;
wire [0:1] mux_tree_tapbuf_size2_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_111_sram;
wire [0:1] mux_tree_tapbuf_size2_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_112_sram;
wire [0:1] mux_tree_tapbuf_size2_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_113_sram;
wire [0:1] mux_tree_tapbuf_size2_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_114_sram;
wire [0:1] mux_tree_tapbuf_size2_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_115_sram;
wire [0:1] mux_tree_tapbuf_size2_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_116_sram;
wire [0:1] mux_tree_tapbuf_size2_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_117_sram;
wire [0:1] mux_tree_tapbuf_size2_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_118_sram;
wire [0:1] mux_tree_tapbuf_size2_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_119_sram;
wire [0:1] mux_tree_tapbuf_size2_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_11_sram;
wire [0:1] mux_tree_tapbuf_size2_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_12_sram;
wire [0:1] mux_tree_tapbuf_size2_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_13_sram;
wire [0:1] mux_tree_tapbuf_size2_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_14_sram;
wire [0:1] mux_tree_tapbuf_size2_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_15_sram;
wire [0:1] mux_tree_tapbuf_size2_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_16_sram;
wire [0:1] mux_tree_tapbuf_size2_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_17_sram;
wire [0:1] mux_tree_tapbuf_size2_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_18_sram;
wire [0:1] mux_tree_tapbuf_size2_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_19_sram;
wire [0:1] mux_tree_tapbuf_size2_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_1_sram;
wire [0:1] mux_tree_tapbuf_size2_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_20_sram;
wire [0:1] mux_tree_tapbuf_size2_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_21_sram;
wire [0:1] mux_tree_tapbuf_size2_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_22_sram;
wire [0:1] mux_tree_tapbuf_size2_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_23_sram;
wire [0:1] mux_tree_tapbuf_size2_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_24_sram;
wire [0:1] mux_tree_tapbuf_size2_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_25_sram;
wire [0:1] mux_tree_tapbuf_size2_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_26_sram;
wire [0:1] mux_tree_tapbuf_size2_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_27_sram;
wire [0:1] mux_tree_tapbuf_size2_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_28_sram;
wire [0:1] mux_tree_tapbuf_size2_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_29_sram;
wire [0:1] mux_tree_tapbuf_size2_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_2_sram;
wire [0:1] mux_tree_tapbuf_size2_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_30_sram;
wire [0:1] mux_tree_tapbuf_size2_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_31_sram;
wire [0:1] mux_tree_tapbuf_size2_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_32_sram;
wire [0:1] mux_tree_tapbuf_size2_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_33_sram;
wire [0:1] mux_tree_tapbuf_size2_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_34_sram;
wire [0:1] mux_tree_tapbuf_size2_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_35_sram;
wire [0:1] mux_tree_tapbuf_size2_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_36_sram;
wire [0:1] mux_tree_tapbuf_size2_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_37_sram;
wire [0:1] mux_tree_tapbuf_size2_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_38_sram;
wire [0:1] mux_tree_tapbuf_size2_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_39_sram;
wire [0:1] mux_tree_tapbuf_size2_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_3_sram;
wire [0:1] mux_tree_tapbuf_size2_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_40_sram;
wire [0:1] mux_tree_tapbuf_size2_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_41_sram;
wire [0:1] mux_tree_tapbuf_size2_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_42_sram;
wire [0:1] mux_tree_tapbuf_size2_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_43_sram;
wire [0:1] mux_tree_tapbuf_size2_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_44_sram;
wire [0:1] mux_tree_tapbuf_size2_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_45_sram;
wire [0:1] mux_tree_tapbuf_size2_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_46_sram;
wire [0:1] mux_tree_tapbuf_size2_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_47_sram;
wire [0:1] mux_tree_tapbuf_size2_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_48_sram;
wire [0:1] mux_tree_tapbuf_size2_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_49_sram;
wire [0:1] mux_tree_tapbuf_size2_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_4_sram;
wire [0:1] mux_tree_tapbuf_size2_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_50_sram;
wire [0:1] mux_tree_tapbuf_size2_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_51_sram;
wire [0:1] mux_tree_tapbuf_size2_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_52_sram;
wire [0:1] mux_tree_tapbuf_size2_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_53_sram;
wire [0:1] mux_tree_tapbuf_size2_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_54_sram;
wire [0:1] mux_tree_tapbuf_size2_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_55_sram;
wire [0:1] mux_tree_tapbuf_size2_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_56_sram;
wire [0:1] mux_tree_tapbuf_size2_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_57_sram;
wire [0:1] mux_tree_tapbuf_size2_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_58_sram;
wire [0:1] mux_tree_tapbuf_size2_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_59_sram;
wire [0:1] mux_tree_tapbuf_size2_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_5_sram;
wire [0:1] mux_tree_tapbuf_size2_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_60_sram;
wire [0:1] mux_tree_tapbuf_size2_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_61_sram;
wire [0:1] mux_tree_tapbuf_size2_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_62_sram;
wire [0:1] mux_tree_tapbuf_size2_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_63_sram;
wire [0:1] mux_tree_tapbuf_size2_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_64_sram;
wire [0:1] mux_tree_tapbuf_size2_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_65_sram;
wire [0:1] mux_tree_tapbuf_size2_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_66_sram;
wire [0:1] mux_tree_tapbuf_size2_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_67_sram;
wire [0:1] mux_tree_tapbuf_size2_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_68_sram;
wire [0:1] mux_tree_tapbuf_size2_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_69_sram;
wire [0:1] mux_tree_tapbuf_size2_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_6_sram;
wire [0:1] mux_tree_tapbuf_size2_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_70_sram;
wire [0:1] mux_tree_tapbuf_size2_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_71_sram;
wire [0:1] mux_tree_tapbuf_size2_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_72_sram;
wire [0:1] mux_tree_tapbuf_size2_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_73_sram;
wire [0:1] mux_tree_tapbuf_size2_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_74_sram;
wire [0:1] mux_tree_tapbuf_size2_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_75_sram;
wire [0:1] mux_tree_tapbuf_size2_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_76_sram;
wire [0:1] mux_tree_tapbuf_size2_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_77_sram;
wire [0:1] mux_tree_tapbuf_size2_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_78_sram;
wire [0:1] mux_tree_tapbuf_size2_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_79_sram;
wire [0:1] mux_tree_tapbuf_size2_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_7_sram;
wire [0:1] mux_tree_tapbuf_size2_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_80_sram;
wire [0:1] mux_tree_tapbuf_size2_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_81_sram;
wire [0:1] mux_tree_tapbuf_size2_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_82_sram;
wire [0:1] mux_tree_tapbuf_size2_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_83_sram;
wire [0:1] mux_tree_tapbuf_size2_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_84_sram;
wire [0:1] mux_tree_tapbuf_size2_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_85_sram;
wire [0:1] mux_tree_tapbuf_size2_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_86_sram;
wire [0:1] mux_tree_tapbuf_size2_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_87_sram;
wire [0:1] mux_tree_tapbuf_size2_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_88_sram;
wire [0:1] mux_tree_tapbuf_size2_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_89_sram;
wire [0:1] mux_tree_tapbuf_size2_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_8_sram;
wire [0:1] mux_tree_tapbuf_size2_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_90_sram;
wire [0:1] mux_tree_tapbuf_size2_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_91_sram;
wire [0:1] mux_tree_tapbuf_size2_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_92_sram;
wire [0:1] mux_tree_tapbuf_size2_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_93_sram;
wire [0:1] mux_tree_tapbuf_size2_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_94_sram;
wire [0:1] mux_tree_tapbuf_size2_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_95_sram;
wire [0:1] mux_tree_tapbuf_size2_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_96_sram;
wire [0:1] mux_tree_tapbuf_size2_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_97_sram;
wire [0:1] mux_tree_tapbuf_size2_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_98_sram;
wire [0:1] mux_tree_tapbuf_size2_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_99_sram;
wire [0:1] mux_tree_tapbuf_size2_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size2_9_sram;
wire [0:1] mux_tree_tapbuf_size2_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size2_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size2_mem_9_ccff_tail;
wire [0:1] mux_tree_tapbuf_size3_0_sram;
wire [0:1] mux_tree_tapbuf_size3_0_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_100_sram;
wire [0:1] mux_tree_tapbuf_size3_100_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_101_sram;
wire [0:1] mux_tree_tapbuf_size3_101_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_102_sram;
wire [0:1] mux_tree_tapbuf_size3_102_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_103_sram;
wire [0:1] mux_tree_tapbuf_size3_103_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_104_sram;
wire [0:1] mux_tree_tapbuf_size3_104_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_105_sram;
wire [0:1] mux_tree_tapbuf_size3_105_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_106_sram;
wire [0:1] mux_tree_tapbuf_size3_106_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_107_sram;
wire [0:1] mux_tree_tapbuf_size3_107_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_108_sram;
wire [0:1] mux_tree_tapbuf_size3_108_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_109_sram;
wire [0:1] mux_tree_tapbuf_size3_109_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_10_sram;
wire [0:1] mux_tree_tapbuf_size3_10_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_110_sram;
wire [0:1] mux_tree_tapbuf_size3_110_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_111_sram;
wire [0:1] mux_tree_tapbuf_size3_111_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_112_sram;
wire [0:1] mux_tree_tapbuf_size3_112_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_113_sram;
wire [0:1] mux_tree_tapbuf_size3_113_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_114_sram;
wire [0:1] mux_tree_tapbuf_size3_114_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_115_sram;
wire [0:1] mux_tree_tapbuf_size3_115_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_116_sram;
wire [0:1] mux_tree_tapbuf_size3_116_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_117_sram;
wire [0:1] mux_tree_tapbuf_size3_117_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_118_sram;
wire [0:1] mux_tree_tapbuf_size3_118_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_119_sram;
wire [0:1] mux_tree_tapbuf_size3_119_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_11_sram;
wire [0:1] mux_tree_tapbuf_size3_11_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_120_sram;
wire [0:1] mux_tree_tapbuf_size3_120_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_121_sram;
wire [0:1] mux_tree_tapbuf_size3_121_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_122_sram;
wire [0:1] mux_tree_tapbuf_size3_122_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_123_sram;
wire [0:1] mux_tree_tapbuf_size3_123_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_124_sram;
wire [0:1] mux_tree_tapbuf_size3_124_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_125_sram;
wire [0:1] mux_tree_tapbuf_size3_125_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_126_sram;
wire [0:1] mux_tree_tapbuf_size3_126_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_127_sram;
wire [0:1] mux_tree_tapbuf_size3_127_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_128_sram;
wire [0:1] mux_tree_tapbuf_size3_128_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_129_sram;
wire [0:1] mux_tree_tapbuf_size3_129_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_12_sram;
wire [0:1] mux_tree_tapbuf_size3_12_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_130_sram;
wire [0:1] mux_tree_tapbuf_size3_130_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_131_sram;
wire [0:1] mux_tree_tapbuf_size3_131_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_132_sram;
wire [0:1] mux_tree_tapbuf_size3_132_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_133_sram;
wire [0:1] mux_tree_tapbuf_size3_133_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_134_sram;
wire [0:1] mux_tree_tapbuf_size3_134_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_135_sram;
wire [0:1] mux_tree_tapbuf_size3_135_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_136_sram;
wire [0:1] mux_tree_tapbuf_size3_136_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_137_sram;
wire [0:1] mux_tree_tapbuf_size3_137_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_138_sram;
wire [0:1] mux_tree_tapbuf_size3_138_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_139_sram;
wire [0:1] mux_tree_tapbuf_size3_139_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_13_sram;
wire [0:1] mux_tree_tapbuf_size3_13_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_140_sram;
wire [0:1] mux_tree_tapbuf_size3_140_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_141_sram;
wire [0:1] mux_tree_tapbuf_size3_141_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_142_sram;
wire [0:1] mux_tree_tapbuf_size3_142_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_143_sram;
wire [0:1] mux_tree_tapbuf_size3_143_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_144_sram;
wire [0:1] mux_tree_tapbuf_size3_144_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_145_sram;
wire [0:1] mux_tree_tapbuf_size3_145_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_146_sram;
wire [0:1] mux_tree_tapbuf_size3_146_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_147_sram;
wire [0:1] mux_tree_tapbuf_size3_147_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_148_sram;
wire [0:1] mux_tree_tapbuf_size3_148_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_149_sram;
wire [0:1] mux_tree_tapbuf_size3_149_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_14_sram;
wire [0:1] mux_tree_tapbuf_size3_14_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_150_sram;
wire [0:1] mux_tree_tapbuf_size3_150_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_151_sram;
wire [0:1] mux_tree_tapbuf_size3_151_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_152_sram;
wire [0:1] mux_tree_tapbuf_size3_152_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_153_sram;
wire [0:1] mux_tree_tapbuf_size3_153_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_154_sram;
wire [0:1] mux_tree_tapbuf_size3_154_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_155_sram;
wire [0:1] mux_tree_tapbuf_size3_155_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_156_sram;
wire [0:1] mux_tree_tapbuf_size3_156_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_157_sram;
wire [0:1] mux_tree_tapbuf_size3_157_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_158_sram;
wire [0:1] mux_tree_tapbuf_size3_158_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_159_sram;
wire [0:1] mux_tree_tapbuf_size3_159_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_15_sram;
wire [0:1] mux_tree_tapbuf_size3_15_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_160_sram;
wire [0:1] mux_tree_tapbuf_size3_160_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_161_sram;
wire [0:1] mux_tree_tapbuf_size3_161_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_162_sram;
wire [0:1] mux_tree_tapbuf_size3_162_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_163_sram;
wire [0:1] mux_tree_tapbuf_size3_163_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_164_sram;
wire [0:1] mux_tree_tapbuf_size3_164_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_165_sram;
wire [0:1] mux_tree_tapbuf_size3_165_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_166_sram;
wire [0:1] mux_tree_tapbuf_size3_166_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_167_sram;
wire [0:1] mux_tree_tapbuf_size3_167_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_168_sram;
wire [0:1] mux_tree_tapbuf_size3_168_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_169_sram;
wire [0:1] mux_tree_tapbuf_size3_169_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_16_sram;
wire [0:1] mux_tree_tapbuf_size3_16_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_170_sram;
wire [0:1] mux_tree_tapbuf_size3_170_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_171_sram;
wire [0:1] mux_tree_tapbuf_size3_171_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_172_sram;
wire [0:1] mux_tree_tapbuf_size3_172_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_173_sram;
wire [0:1] mux_tree_tapbuf_size3_173_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_174_sram;
wire [0:1] mux_tree_tapbuf_size3_174_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_175_sram;
wire [0:1] mux_tree_tapbuf_size3_175_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_176_sram;
wire [0:1] mux_tree_tapbuf_size3_176_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_177_sram;
wire [0:1] mux_tree_tapbuf_size3_177_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_178_sram;
wire [0:1] mux_tree_tapbuf_size3_178_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_179_sram;
wire [0:1] mux_tree_tapbuf_size3_179_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_17_sram;
wire [0:1] mux_tree_tapbuf_size3_17_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_180_sram;
wire [0:1] mux_tree_tapbuf_size3_180_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_181_sram;
wire [0:1] mux_tree_tapbuf_size3_181_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_182_sram;
wire [0:1] mux_tree_tapbuf_size3_182_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_183_sram;
wire [0:1] mux_tree_tapbuf_size3_183_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_184_sram;
wire [0:1] mux_tree_tapbuf_size3_184_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_185_sram;
wire [0:1] mux_tree_tapbuf_size3_185_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_186_sram;
wire [0:1] mux_tree_tapbuf_size3_186_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_187_sram;
wire [0:1] mux_tree_tapbuf_size3_187_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_188_sram;
wire [0:1] mux_tree_tapbuf_size3_188_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_189_sram;
wire [0:1] mux_tree_tapbuf_size3_189_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_18_sram;
wire [0:1] mux_tree_tapbuf_size3_18_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_190_sram;
wire [0:1] mux_tree_tapbuf_size3_190_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_191_sram;
wire [0:1] mux_tree_tapbuf_size3_191_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_192_sram;
wire [0:1] mux_tree_tapbuf_size3_192_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_193_sram;
wire [0:1] mux_tree_tapbuf_size3_193_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_194_sram;
wire [0:1] mux_tree_tapbuf_size3_194_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_195_sram;
wire [0:1] mux_tree_tapbuf_size3_195_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_196_sram;
wire [0:1] mux_tree_tapbuf_size3_196_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_197_sram;
wire [0:1] mux_tree_tapbuf_size3_197_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_198_sram;
wire [0:1] mux_tree_tapbuf_size3_198_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_199_sram;
wire [0:1] mux_tree_tapbuf_size3_199_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_19_sram;
wire [0:1] mux_tree_tapbuf_size3_19_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_1_sram;
wire [0:1] mux_tree_tapbuf_size3_1_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_200_sram;
wire [0:1] mux_tree_tapbuf_size3_200_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_201_sram;
wire [0:1] mux_tree_tapbuf_size3_201_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_202_sram;
wire [0:1] mux_tree_tapbuf_size3_202_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_203_sram;
wire [0:1] mux_tree_tapbuf_size3_203_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_204_sram;
wire [0:1] mux_tree_tapbuf_size3_204_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_205_sram;
wire [0:1] mux_tree_tapbuf_size3_205_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_206_sram;
wire [0:1] mux_tree_tapbuf_size3_206_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_207_sram;
wire [0:1] mux_tree_tapbuf_size3_207_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_208_sram;
wire [0:1] mux_tree_tapbuf_size3_208_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_209_sram;
wire [0:1] mux_tree_tapbuf_size3_209_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_20_sram;
wire [0:1] mux_tree_tapbuf_size3_20_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_210_sram;
wire [0:1] mux_tree_tapbuf_size3_210_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_211_sram;
wire [0:1] mux_tree_tapbuf_size3_211_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_212_sram;
wire [0:1] mux_tree_tapbuf_size3_212_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_213_sram;
wire [0:1] mux_tree_tapbuf_size3_213_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_214_sram;
wire [0:1] mux_tree_tapbuf_size3_214_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_215_sram;
wire [0:1] mux_tree_tapbuf_size3_215_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_216_sram;
wire [0:1] mux_tree_tapbuf_size3_216_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_217_sram;
wire [0:1] mux_tree_tapbuf_size3_217_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_218_sram;
wire [0:1] mux_tree_tapbuf_size3_218_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_219_sram;
wire [0:1] mux_tree_tapbuf_size3_219_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_21_sram;
wire [0:1] mux_tree_tapbuf_size3_21_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_220_sram;
wire [0:1] mux_tree_tapbuf_size3_220_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_221_sram;
wire [0:1] mux_tree_tapbuf_size3_221_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_222_sram;
wire [0:1] mux_tree_tapbuf_size3_222_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_223_sram;
wire [0:1] mux_tree_tapbuf_size3_223_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_224_sram;
wire [0:1] mux_tree_tapbuf_size3_224_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_225_sram;
wire [0:1] mux_tree_tapbuf_size3_225_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_226_sram;
wire [0:1] mux_tree_tapbuf_size3_226_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_227_sram;
wire [0:1] mux_tree_tapbuf_size3_227_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_228_sram;
wire [0:1] mux_tree_tapbuf_size3_228_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_229_sram;
wire [0:1] mux_tree_tapbuf_size3_229_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_22_sram;
wire [0:1] mux_tree_tapbuf_size3_22_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_230_sram;
wire [0:1] mux_tree_tapbuf_size3_230_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_231_sram;
wire [0:1] mux_tree_tapbuf_size3_231_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_232_sram;
wire [0:1] mux_tree_tapbuf_size3_232_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_233_sram;
wire [0:1] mux_tree_tapbuf_size3_233_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_234_sram;
wire [0:1] mux_tree_tapbuf_size3_234_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_235_sram;
wire [0:1] mux_tree_tapbuf_size3_235_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_236_sram;
wire [0:1] mux_tree_tapbuf_size3_236_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_237_sram;
wire [0:1] mux_tree_tapbuf_size3_237_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_238_sram;
wire [0:1] mux_tree_tapbuf_size3_238_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_239_sram;
wire [0:1] mux_tree_tapbuf_size3_239_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_23_sram;
wire [0:1] mux_tree_tapbuf_size3_23_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_240_sram;
wire [0:1] mux_tree_tapbuf_size3_240_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_241_sram;
wire [0:1] mux_tree_tapbuf_size3_241_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_242_sram;
wire [0:1] mux_tree_tapbuf_size3_242_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_243_sram;
wire [0:1] mux_tree_tapbuf_size3_243_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_244_sram;
wire [0:1] mux_tree_tapbuf_size3_244_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_245_sram;
wire [0:1] mux_tree_tapbuf_size3_245_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_246_sram;
wire [0:1] mux_tree_tapbuf_size3_246_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_247_sram;
wire [0:1] mux_tree_tapbuf_size3_247_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_248_sram;
wire [0:1] mux_tree_tapbuf_size3_248_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_249_sram;
wire [0:1] mux_tree_tapbuf_size3_249_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_24_sram;
wire [0:1] mux_tree_tapbuf_size3_24_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_250_sram;
wire [0:1] mux_tree_tapbuf_size3_250_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_251_sram;
wire [0:1] mux_tree_tapbuf_size3_251_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_252_sram;
wire [0:1] mux_tree_tapbuf_size3_252_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_253_sram;
wire [0:1] mux_tree_tapbuf_size3_253_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_254_sram;
wire [0:1] mux_tree_tapbuf_size3_254_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_255_sram;
wire [0:1] mux_tree_tapbuf_size3_255_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_256_sram;
wire [0:1] mux_tree_tapbuf_size3_256_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_257_sram;
wire [0:1] mux_tree_tapbuf_size3_257_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_258_sram;
wire [0:1] mux_tree_tapbuf_size3_258_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_259_sram;
wire [0:1] mux_tree_tapbuf_size3_259_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_25_sram;
wire [0:1] mux_tree_tapbuf_size3_25_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_260_sram;
wire [0:1] mux_tree_tapbuf_size3_260_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_261_sram;
wire [0:1] mux_tree_tapbuf_size3_261_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_262_sram;
wire [0:1] mux_tree_tapbuf_size3_262_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_263_sram;
wire [0:1] mux_tree_tapbuf_size3_263_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_264_sram;
wire [0:1] mux_tree_tapbuf_size3_264_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_265_sram;
wire [0:1] mux_tree_tapbuf_size3_265_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_266_sram;
wire [0:1] mux_tree_tapbuf_size3_266_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_267_sram;
wire [0:1] mux_tree_tapbuf_size3_267_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_268_sram;
wire [0:1] mux_tree_tapbuf_size3_268_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_269_sram;
wire [0:1] mux_tree_tapbuf_size3_269_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_26_sram;
wire [0:1] mux_tree_tapbuf_size3_26_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_270_sram;
wire [0:1] mux_tree_tapbuf_size3_270_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_271_sram;
wire [0:1] mux_tree_tapbuf_size3_271_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_272_sram;
wire [0:1] mux_tree_tapbuf_size3_272_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_273_sram;
wire [0:1] mux_tree_tapbuf_size3_273_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_274_sram;
wire [0:1] mux_tree_tapbuf_size3_274_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_275_sram;
wire [0:1] mux_tree_tapbuf_size3_275_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_276_sram;
wire [0:1] mux_tree_tapbuf_size3_276_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_277_sram;
wire [0:1] mux_tree_tapbuf_size3_277_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_278_sram;
wire [0:1] mux_tree_tapbuf_size3_278_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_279_sram;
wire [0:1] mux_tree_tapbuf_size3_279_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_27_sram;
wire [0:1] mux_tree_tapbuf_size3_27_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_280_sram;
wire [0:1] mux_tree_tapbuf_size3_280_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_281_sram;
wire [0:1] mux_tree_tapbuf_size3_281_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_282_sram;
wire [0:1] mux_tree_tapbuf_size3_282_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_283_sram;
wire [0:1] mux_tree_tapbuf_size3_283_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_284_sram;
wire [0:1] mux_tree_tapbuf_size3_284_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_285_sram;
wire [0:1] mux_tree_tapbuf_size3_285_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_286_sram;
wire [0:1] mux_tree_tapbuf_size3_286_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_287_sram;
wire [0:1] mux_tree_tapbuf_size3_287_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_288_sram;
wire [0:1] mux_tree_tapbuf_size3_288_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_289_sram;
wire [0:1] mux_tree_tapbuf_size3_289_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_28_sram;
wire [0:1] mux_tree_tapbuf_size3_28_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_290_sram;
wire [0:1] mux_tree_tapbuf_size3_290_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_291_sram;
wire [0:1] mux_tree_tapbuf_size3_291_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_292_sram;
wire [0:1] mux_tree_tapbuf_size3_292_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_293_sram;
wire [0:1] mux_tree_tapbuf_size3_293_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_294_sram;
wire [0:1] mux_tree_tapbuf_size3_294_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_295_sram;
wire [0:1] mux_tree_tapbuf_size3_295_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_296_sram;
wire [0:1] mux_tree_tapbuf_size3_296_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_297_sram;
wire [0:1] mux_tree_tapbuf_size3_297_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_298_sram;
wire [0:1] mux_tree_tapbuf_size3_298_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_299_sram;
wire [0:1] mux_tree_tapbuf_size3_299_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_29_sram;
wire [0:1] mux_tree_tapbuf_size3_29_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_2_sram;
wire [0:1] mux_tree_tapbuf_size3_2_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_300_sram;
wire [0:1] mux_tree_tapbuf_size3_300_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_301_sram;
wire [0:1] mux_tree_tapbuf_size3_301_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_302_sram;
wire [0:1] mux_tree_tapbuf_size3_302_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_303_sram;
wire [0:1] mux_tree_tapbuf_size3_303_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_304_sram;
wire [0:1] mux_tree_tapbuf_size3_304_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_305_sram;
wire [0:1] mux_tree_tapbuf_size3_305_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_306_sram;
wire [0:1] mux_tree_tapbuf_size3_306_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_307_sram;
wire [0:1] mux_tree_tapbuf_size3_307_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_308_sram;
wire [0:1] mux_tree_tapbuf_size3_308_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_309_sram;
wire [0:1] mux_tree_tapbuf_size3_309_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_30_sram;
wire [0:1] mux_tree_tapbuf_size3_30_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_310_sram;
wire [0:1] mux_tree_tapbuf_size3_310_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_311_sram;
wire [0:1] mux_tree_tapbuf_size3_311_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_312_sram;
wire [0:1] mux_tree_tapbuf_size3_312_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_313_sram;
wire [0:1] mux_tree_tapbuf_size3_313_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_314_sram;
wire [0:1] mux_tree_tapbuf_size3_314_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_315_sram;
wire [0:1] mux_tree_tapbuf_size3_315_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_316_sram;
wire [0:1] mux_tree_tapbuf_size3_316_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_317_sram;
wire [0:1] mux_tree_tapbuf_size3_317_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_318_sram;
wire [0:1] mux_tree_tapbuf_size3_318_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_319_sram;
wire [0:1] mux_tree_tapbuf_size3_319_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_31_sram;
wire [0:1] mux_tree_tapbuf_size3_31_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_320_sram;
wire [0:1] mux_tree_tapbuf_size3_320_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_321_sram;
wire [0:1] mux_tree_tapbuf_size3_321_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_322_sram;
wire [0:1] mux_tree_tapbuf_size3_322_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_323_sram;
wire [0:1] mux_tree_tapbuf_size3_323_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_324_sram;
wire [0:1] mux_tree_tapbuf_size3_324_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_325_sram;
wire [0:1] mux_tree_tapbuf_size3_325_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_326_sram;
wire [0:1] mux_tree_tapbuf_size3_326_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_327_sram;
wire [0:1] mux_tree_tapbuf_size3_327_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_328_sram;
wire [0:1] mux_tree_tapbuf_size3_328_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_329_sram;
wire [0:1] mux_tree_tapbuf_size3_329_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_32_sram;
wire [0:1] mux_tree_tapbuf_size3_32_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_330_sram;
wire [0:1] mux_tree_tapbuf_size3_330_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_331_sram;
wire [0:1] mux_tree_tapbuf_size3_331_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_332_sram;
wire [0:1] mux_tree_tapbuf_size3_332_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_333_sram;
wire [0:1] mux_tree_tapbuf_size3_333_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_334_sram;
wire [0:1] mux_tree_tapbuf_size3_334_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_335_sram;
wire [0:1] mux_tree_tapbuf_size3_335_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_336_sram;
wire [0:1] mux_tree_tapbuf_size3_336_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_337_sram;
wire [0:1] mux_tree_tapbuf_size3_337_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_338_sram;
wire [0:1] mux_tree_tapbuf_size3_338_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_339_sram;
wire [0:1] mux_tree_tapbuf_size3_339_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_33_sram;
wire [0:1] mux_tree_tapbuf_size3_33_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_340_sram;
wire [0:1] mux_tree_tapbuf_size3_340_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_341_sram;
wire [0:1] mux_tree_tapbuf_size3_341_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_342_sram;
wire [0:1] mux_tree_tapbuf_size3_342_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_343_sram;
wire [0:1] mux_tree_tapbuf_size3_343_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_344_sram;
wire [0:1] mux_tree_tapbuf_size3_344_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_345_sram;
wire [0:1] mux_tree_tapbuf_size3_345_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_346_sram;
wire [0:1] mux_tree_tapbuf_size3_346_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_347_sram;
wire [0:1] mux_tree_tapbuf_size3_347_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_348_sram;
wire [0:1] mux_tree_tapbuf_size3_348_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_349_sram;
wire [0:1] mux_tree_tapbuf_size3_349_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_34_sram;
wire [0:1] mux_tree_tapbuf_size3_34_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_350_sram;
wire [0:1] mux_tree_tapbuf_size3_350_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_351_sram;
wire [0:1] mux_tree_tapbuf_size3_351_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_352_sram;
wire [0:1] mux_tree_tapbuf_size3_352_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_353_sram;
wire [0:1] mux_tree_tapbuf_size3_353_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_354_sram;
wire [0:1] mux_tree_tapbuf_size3_354_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_355_sram;
wire [0:1] mux_tree_tapbuf_size3_355_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_356_sram;
wire [0:1] mux_tree_tapbuf_size3_356_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_357_sram;
wire [0:1] mux_tree_tapbuf_size3_357_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_358_sram;
wire [0:1] mux_tree_tapbuf_size3_358_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_359_sram;
wire [0:1] mux_tree_tapbuf_size3_359_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_35_sram;
wire [0:1] mux_tree_tapbuf_size3_35_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_360_sram;
wire [0:1] mux_tree_tapbuf_size3_360_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_361_sram;
wire [0:1] mux_tree_tapbuf_size3_361_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_362_sram;
wire [0:1] mux_tree_tapbuf_size3_362_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_363_sram;
wire [0:1] mux_tree_tapbuf_size3_363_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_364_sram;
wire [0:1] mux_tree_tapbuf_size3_364_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_365_sram;
wire [0:1] mux_tree_tapbuf_size3_365_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_366_sram;
wire [0:1] mux_tree_tapbuf_size3_366_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_367_sram;
wire [0:1] mux_tree_tapbuf_size3_367_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_368_sram;
wire [0:1] mux_tree_tapbuf_size3_368_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_369_sram;
wire [0:1] mux_tree_tapbuf_size3_369_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_36_sram;
wire [0:1] mux_tree_tapbuf_size3_36_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_370_sram;
wire [0:1] mux_tree_tapbuf_size3_370_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_371_sram;
wire [0:1] mux_tree_tapbuf_size3_371_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_372_sram;
wire [0:1] mux_tree_tapbuf_size3_372_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_373_sram;
wire [0:1] mux_tree_tapbuf_size3_373_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_374_sram;
wire [0:1] mux_tree_tapbuf_size3_374_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_375_sram;
wire [0:1] mux_tree_tapbuf_size3_375_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_376_sram;
wire [0:1] mux_tree_tapbuf_size3_376_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_377_sram;
wire [0:1] mux_tree_tapbuf_size3_377_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_378_sram;
wire [0:1] mux_tree_tapbuf_size3_378_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_379_sram;
wire [0:1] mux_tree_tapbuf_size3_379_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_37_sram;
wire [0:1] mux_tree_tapbuf_size3_37_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_380_sram;
wire [0:1] mux_tree_tapbuf_size3_380_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_381_sram;
wire [0:1] mux_tree_tapbuf_size3_381_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_382_sram;
wire [0:1] mux_tree_tapbuf_size3_382_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_383_sram;
wire [0:1] mux_tree_tapbuf_size3_383_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_384_sram;
wire [0:1] mux_tree_tapbuf_size3_384_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_385_sram;
wire [0:1] mux_tree_tapbuf_size3_385_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_386_sram;
wire [0:1] mux_tree_tapbuf_size3_386_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_387_sram;
wire [0:1] mux_tree_tapbuf_size3_387_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_388_sram;
wire [0:1] mux_tree_tapbuf_size3_388_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_389_sram;
wire [0:1] mux_tree_tapbuf_size3_389_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_38_sram;
wire [0:1] mux_tree_tapbuf_size3_38_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_390_sram;
wire [0:1] mux_tree_tapbuf_size3_390_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_391_sram;
wire [0:1] mux_tree_tapbuf_size3_391_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_392_sram;
wire [0:1] mux_tree_tapbuf_size3_392_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_393_sram;
wire [0:1] mux_tree_tapbuf_size3_393_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_394_sram;
wire [0:1] mux_tree_tapbuf_size3_394_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_395_sram;
wire [0:1] mux_tree_tapbuf_size3_395_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_396_sram;
wire [0:1] mux_tree_tapbuf_size3_396_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_397_sram;
wire [0:1] mux_tree_tapbuf_size3_397_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_398_sram;
wire [0:1] mux_tree_tapbuf_size3_398_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_399_sram;
wire [0:1] mux_tree_tapbuf_size3_399_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_39_sram;
wire [0:1] mux_tree_tapbuf_size3_39_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_3_sram;
wire [0:1] mux_tree_tapbuf_size3_3_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_400_sram;
wire [0:1] mux_tree_tapbuf_size3_400_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_401_sram;
wire [0:1] mux_tree_tapbuf_size3_401_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_402_sram;
wire [0:1] mux_tree_tapbuf_size3_402_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_403_sram;
wire [0:1] mux_tree_tapbuf_size3_403_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_404_sram;
wire [0:1] mux_tree_tapbuf_size3_404_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_405_sram;
wire [0:1] mux_tree_tapbuf_size3_405_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_406_sram;
wire [0:1] mux_tree_tapbuf_size3_406_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_407_sram;
wire [0:1] mux_tree_tapbuf_size3_407_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_408_sram;
wire [0:1] mux_tree_tapbuf_size3_408_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_409_sram;
wire [0:1] mux_tree_tapbuf_size3_409_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_40_sram;
wire [0:1] mux_tree_tapbuf_size3_40_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_410_sram;
wire [0:1] mux_tree_tapbuf_size3_410_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_411_sram;
wire [0:1] mux_tree_tapbuf_size3_411_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_412_sram;
wire [0:1] mux_tree_tapbuf_size3_412_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_413_sram;
wire [0:1] mux_tree_tapbuf_size3_413_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_414_sram;
wire [0:1] mux_tree_tapbuf_size3_414_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_415_sram;
wire [0:1] mux_tree_tapbuf_size3_415_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_416_sram;
wire [0:1] mux_tree_tapbuf_size3_416_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_417_sram;
wire [0:1] mux_tree_tapbuf_size3_417_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_418_sram;
wire [0:1] mux_tree_tapbuf_size3_418_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_419_sram;
wire [0:1] mux_tree_tapbuf_size3_419_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_41_sram;
wire [0:1] mux_tree_tapbuf_size3_41_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_420_sram;
wire [0:1] mux_tree_tapbuf_size3_420_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_421_sram;
wire [0:1] mux_tree_tapbuf_size3_421_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_422_sram;
wire [0:1] mux_tree_tapbuf_size3_422_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_423_sram;
wire [0:1] mux_tree_tapbuf_size3_423_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_424_sram;
wire [0:1] mux_tree_tapbuf_size3_424_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_425_sram;
wire [0:1] mux_tree_tapbuf_size3_425_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_426_sram;
wire [0:1] mux_tree_tapbuf_size3_426_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_427_sram;
wire [0:1] mux_tree_tapbuf_size3_427_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_428_sram;
wire [0:1] mux_tree_tapbuf_size3_428_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_429_sram;
wire [0:1] mux_tree_tapbuf_size3_429_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_42_sram;
wire [0:1] mux_tree_tapbuf_size3_42_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_430_sram;
wire [0:1] mux_tree_tapbuf_size3_430_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_431_sram;
wire [0:1] mux_tree_tapbuf_size3_431_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_432_sram;
wire [0:1] mux_tree_tapbuf_size3_432_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_433_sram;
wire [0:1] mux_tree_tapbuf_size3_433_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_434_sram;
wire [0:1] mux_tree_tapbuf_size3_434_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_435_sram;
wire [0:1] mux_tree_tapbuf_size3_435_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_436_sram;
wire [0:1] mux_tree_tapbuf_size3_436_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_437_sram;
wire [0:1] mux_tree_tapbuf_size3_437_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_438_sram;
wire [0:1] mux_tree_tapbuf_size3_438_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_439_sram;
wire [0:1] mux_tree_tapbuf_size3_439_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_43_sram;
wire [0:1] mux_tree_tapbuf_size3_43_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_440_sram;
wire [0:1] mux_tree_tapbuf_size3_440_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_441_sram;
wire [0:1] mux_tree_tapbuf_size3_441_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_442_sram;
wire [0:1] mux_tree_tapbuf_size3_442_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_443_sram;
wire [0:1] mux_tree_tapbuf_size3_443_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_444_sram;
wire [0:1] mux_tree_tapbuf_size3_444_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_445_sram;
wire [0:1] mux_tree_tapbuf_size3_445_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_44_sram;
wire [0:1] mux_tree_tapbuf_size3_44_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_45_sram;
wire [0:1] mux_tree_tapbuf_size3_45_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_46_sram;
wire [0:1] mux_tree_tapbuf_size3_46_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_47_sram;
wire [0:1] mux_tree_tapbuf_size3_47_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_48_sram;
wire [0:1] mux_tree_tapbuf_size3_48_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_49_sram;
wire [0:1] mux_tree_tapbuf_size3_49_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_4_sram;
wire [0:1] mux_tree_tapbuf_size3_4_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_50_sram;
wire [0:1] mux_tree_tapbuf_size3_50_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_51_sram;
wire [0:1] mux_tree_tapbuf_size3_51_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_52_sram;
wire [0:1] mux_tree_tapbuf_size3_52_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_53_sram;
wire [0:1] mux_tree_tapbuf_size3_53_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_54_sram;
wire [0:1] mux_tree_tapbuf_size3_54_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_55_sram;
wire [0:1] mux_tree_tapbuf_size3_55_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_56_sram;
wire [0:1] mux_tree_tapbuf_size3_56_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_57_sram;
wire [0:1] mux_tree_tapbuf_size3_57_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_58_sram;
wire [0:1] mux_tree_tapbuf_size3_58_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_59_sram;
wire [0:1] mux_tree_tapbuf_size3_59_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_5_sram;
wire [0:1] mux_tree_tapbuf_size3_5_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_60_sram;
wire [0:1] mux_tree_tapbuf_size3_60_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_61_sram;
wire [0:1] mux_tree_tapbuf_size3_61_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_62_sram;
wire [0:1] mux_tree_tapbuf_size3_62_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_63_sram;
wire [0:1] mux_tree_tapbuf_size3_63_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_64_sram;
wire [0:1] mux_tree_tapbuf_size3_64_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_65_sram;
wire [0:1] mux_tree_tapbuf_size3_65_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_66_sram;
wire [0:1] mux_tree_tapbuf_size3_66_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_67_sram;
wire [0:1] mux_tree_tapbuf_size3_67_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_68_sram;
wire [0:1] mux_tree_tapbuf_size3_68_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_69_sram;
wire [0:1] mux_tree_tapbuf_size3_69_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_6_sram;
wire [0:1] mux_tree_tapbuf_size3_6_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_70_sram;
wire [0:1] mux_tree_tapbuf_size3_70_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_71_sram;
wire [0:1] mux_tree_tapbuf_size3_71_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_72_sram;
wire [0:1] mux_tree_tapbuf_size3_72_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_73_sram;
wire [0:1] mux_tree_tapbuf_size3_73_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_74_sram;
wire [0:1] mux_tree_tapbuf_size3_74_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_75_sram;
wire [0:1] mux_tree_tapbuf_size3_75_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_76_sram;
wire [0:1] mux_tree_tapbuf_size3_76_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_77_sram;
wire [0:1] mux_tree_tapbuf_size3_77_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_78_sram;
wire [0:1] mux_tree_tapbuf_size3_78_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_79_sram;
wire [0:1] mux_tree_tapbuf_size3_79_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_7_sram;
wire [0:1] mux_tree_tapbuf_size3_7_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_80_sram;
wire [0:1] mux_tree_tapbuf_size3_80_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_81_sram;
wire [0:1] mux_tree_tapbuf_size3_81_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_82_sram;
wire [0:1] mux_tree_tapbuf_size3_82_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_83_sram;
wire [0:1] mux_tree_tapbuf_size3_83_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_84_sram;
wire [0:1] mux_tree_tapbuf_size3_84_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_85_sram;
wire [0:1] mux_tree_tapbuf_size3_85_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_86_sram;
wire [0:1] mux_tree_tapbuf_size3_86_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_87_sram;
wire [0:1] mux_tree_tapbuf_size3_87_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_88_sram;
wire [0:1] mux_tree_tapbuf_size3_88_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_89_sram;
wire [0:1] mux_tree_tapbuf_size3_89_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_8_sram;
wire [0:1] mux_tree_tapbuf_size3_8_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_90_sram;
wire [0:1] mux_tree_tapbuf_size3_90_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_91_sram;
wire [0:1] mux_tree_tapbuf_size3_91_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_92_sram;
wire [0:1] mux_tree_tapbuf_size3_92_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_93_sram;
wire [0:1] mux_tree_tapbuf_size3_93_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_94_sram;
wire [0:1] mux_tree_tapbuf_size3_94_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_95_sram;
wire [0:1] mux_tree_tapbuf_size3_95_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_96_sram;
wire [0:1] mux_tree_tapbuf_size3_96_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_97_sram;
wire [0:1] mux_tree_tapbuf_size3_97_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_98_sram;
wire [0:1] mux_tree_tapbuf_size3_98_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_99_sram;
wire [0:1] mux_tree_tapbuf_size3_99_sram_inv;
wire [0:1] mux_tree_tapbuf_size3_9_sram;
wire [0:1] mux_tree_tapbuf_size3_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size3_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_100_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_101_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_102_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_103_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_104_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_105_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_106_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_107_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_108_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_109_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_110_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_111_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_112_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_113_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_114_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_115_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_116_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_117_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_118_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_119_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_120_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_121_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_122_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_123_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_124_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_125_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_126_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_127_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_128_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_129_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_130_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_131_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_132_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_133_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_134_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_135_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_136_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_137_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_138_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_139_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_140_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_141_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_142_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_143_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_144_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_145_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_146_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_147_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_148_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_149_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_150_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_151_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_152_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_153_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_154_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_155_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_156_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_157_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_158_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_159_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_160_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_161_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_162_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_163_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_164_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_165_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_166_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_167_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_168_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_169_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_170_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_171_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_172_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_173_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_174_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_175_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_176_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_177_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_178_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_179_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_180_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_181_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_182_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_183_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_184_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_185_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_186_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_187_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_188_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_189_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_190_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_191_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_192_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_193_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_194_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_195_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_196_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_197_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_198_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_199_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_200_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_201_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_202_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_203_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_204_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_205_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_206_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_207_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_208_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_209_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_210_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_211_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_212_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_213_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_214_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_215_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_216_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_217_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_218_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_219_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_220_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_221_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_222_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_223_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_224_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_225_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_226_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_227_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_228_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_229_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_230_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_231_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_232_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_233_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_234_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_235_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_236_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_237_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_238_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_239_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_240_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_241_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_242_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_243_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_244_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_245_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_246_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_247_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_248_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_249_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_250_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_251_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_252_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_253_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_254_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_255_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_256_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_257_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_258_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_259_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_260_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_261_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_262_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_263_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_264_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_265_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_266_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_267_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_268_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_269_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_270_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_271_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_272_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_273_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_274_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_275_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_276_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_277_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_278_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_279_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_280_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_281_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_282_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_283_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_284_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_285_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_286_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_287_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_288_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_289_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_290_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_291_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_292_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_293_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_294_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_295_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_296_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_297_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_298_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_299_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_300_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_301_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_302_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_303_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_304_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_305_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_306_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_307_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_308_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_309_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_310_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_311_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_312_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_313_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_314_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_315_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_316_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_317_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_318_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_319_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_320_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_321_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_322_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_323_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_324_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_325_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_326_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_327_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_328_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_329_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_330_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_331_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_332_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_333_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_334_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_335_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_336_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_337_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_338_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_339_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_340_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_341_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_342_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_343_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_344_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_345_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_346_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_347_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_348_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_349_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_350_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_351_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_352_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_353_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_354_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_355_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_356_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_357_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_358_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_359_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_360_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_361_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_362_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_363_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_364_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_365_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_366_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_367_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_368_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_369_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_370_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_371_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_372_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_373_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_374_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_375_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_376_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_377_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_378_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_379_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_37_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_380_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_381_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_382_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_383_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_384_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_385_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_386_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_387_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_388_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_389_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_38_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_390_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_391_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_392_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_393_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_394_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_395_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_396_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_397_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_398_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_399_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_39_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_400_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_401_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_402_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_403_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_404_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_405_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_406_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_407_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_408_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_409_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_40_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_410_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_411_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_412_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_413_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_414_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_415_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_416_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_417_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_418_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_419_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_41_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_420_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_421_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_422_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_423_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_424_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_425_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_426_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_427_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_428_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_429_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_42_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_430_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_431_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_432_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_433_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_434_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_435_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_436_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_437_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_438_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_439_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_43_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_440_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_441_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_442_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_443_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_444_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_44_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_45_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_46_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_47_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_48_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_49_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_50_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_51_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_52_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_53_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_54_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_55_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_56_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_57_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_58_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_59_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_60_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_61_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_62_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_63_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_64_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_65_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_66_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_67_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_68_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_69_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_70_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_71_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_72_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_73_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_74_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_75_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_76_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_77_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_78_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_79_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_80_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_81_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_82_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_83_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_84_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_85_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_86_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_87_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_88_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_89_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_90_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_91_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_92_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_93_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_94_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_95_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_96_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_97_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_98_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_99_ccff_tail;
wire [0:0] mux_tree_tapbuf_size3_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size4_0_sram;
wire [0:2] mux_tree_tapbuf_size4_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_1_sram;
wire [0:2] mux_tree_tapbuf_size4_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_2_sram;
wire [0:2] mux_tree_tapbuf_size4_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size4_3_sram;
wire [0:2] mux_tree_tapbuf_size4_3_sram_inv;
wire [0:0] mux_tree_tapbuf_size4_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size4_mem_3_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size4 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[1]}),
		.sram(mux_tree_tapbuf_size4_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_0_sram_inv[0:2]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size4 mux_top_track_18 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[10]}),
		.sram(mux_tree_tapbuf_size4_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_1_sram_inv[0:2]),
		.out(chany_top_out[9]));

	mux_tree_tapbuf_size4 mux_right_track_0 (
		.in({chany_top_in[284], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_2_sram_inv[0:2]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size4 mux_right_track_18 (
		.in({chany_top_in[8], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size4_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size4_3_sram_inv[0:2]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size4_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_0_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_top_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_1_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_222_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_2_sram_inv[0:2]));

	mux_tree_tapbuf_size4_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_230_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size4_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size4_3_sram_inv[0:2]));

	mux_tree_tapbuf_size3 mux_top_track_2 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[2]}),
		.sram(mux_tree_tapbuf_size3_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_0_sram_inv[0:1]),
		.out(chany_top_out[1]));

	mux_tree_tapbuf_size3 mux_top_track_4 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[3]}),
		.sram(mux_tree_tapbuf_size3_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_1_sram_inv[0:1]),
		.out(chany_top_out[2]));

	mux_tree_tapbuf_size3 mux_top_track_6 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[4]}),
		.sram(mux_tree_tapbuf_size3_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_2_sram_inv[0:1]),
		.out(chany_top_out[3]));

	mux_tree_tapbuf_size3 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[5]}),
		.sram(mux_tree_tapbuf_size3_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_3_sram_inv[0:1]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size3 mux_top_track_10 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[6]}),
		.sram(mux_tree_tapbuf_size3_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_4_sram_inv[0:1]),
		.out(chany_top_out[5]));

	mux_tree_tapbuf_size3 mux_top_track_12 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[7]}),
		.sram(mux_tree_tapbuf_size3_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_5_sram_inv[0:1]),
		.out(chany_top_out[6]));

	mux_tree_tapbuf_size3 mux_top_track_14 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[8]}),
		.sram(mux_tree_tapbuf_size3_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_6_sram_inv[0:1]),
		.out(chany_top_out[7]));

	mux_tree_tapbuf_size3 mux_top_track_16 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[9]}),
		.sram(mux_tree_tapbuf_size3_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_7_sram_inv[0:1]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size3 mux_top_track_20 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[11]}),
		.sram(mux_tree_tapbuf_size3_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_8_sram_inv[0:1]),
		.out(chany_top_out[10]));

	mux_tree_tapbuf_size3 mux_top_track_22 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[12]}),
		.sram(mux_tree_tapbuf_size3_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_9_sram_inv[0:1]),
		.out(chany_top_out[11]));

	mux_tree_tapbuf_size3 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[13]}),
		.sram(mux_tree_tapbuf_size3_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_10_sram_inv[0:1]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size3 mux_top_track_26 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[14]}),
		.sram(mux_tree_tapbuf_size3_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_11_sram_inv[0:1]),
		.out(chany_top_out[13]));

	mux_tree_tapbuf_size3 mux_top_track_28 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[15]}),
		.sram(mux_tree_tapbuf_size3_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_12_sram_inv[0:1]),
		.out(chany_top_out[14]));

	mux_tree_tapbuf_size3 mux_top_track_30 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[16]}),
		.sram(mux_tree_tapbuf_size3_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_13_sram_inv[0:1]),
		.out(chany_top_out[15]));

	mux_tree_tapbuf_size3 mux_top_track_36 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[19]}),
		.sram(mux_tree_tapbuf_size3_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_14_sram_inv[0:1]),
		.out(chany_top_out[18]));

	mux_tree_tapbuf_size3 mux_top_track_38 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[20]}),
		.sram(mux_tree_tapbuf_size3_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_15_sram_inv[0:1]),
		.out(chany_top_out[19]));

	mux_tree_tapbuf_size3 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[21]}),
		.sram(mux_tree_tapbuf_size3_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_16_sram_inv[0:1]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size3 mux_top_track_42 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[22]}),
		.sram(mux_tree_tapbuf_size3_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_17_sram_inv[0:1]),
		.out(chany_top_out[21]));

	mux_tree_tapbuf_size3 mux_top_track_44 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[23]}),
		.sram(mux_tree_tapbuf_size3_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_18_sram_inv[0:1]),
		.out(chany_top_out[22]));

	mux_tree_tapbuf_size3 mux_top_track_46 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[24]}),
		.sram(mux_tree_tapbuf_size3_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_19_sram_inv[0:1]),
		.out(chany_top_out[23]));

	mux_tree_tapbuf_size3 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[25]}),
		.sram(mux_tree_tapbuf_size3_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_20_sram_inv[0:1]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size3 mux_top_track_54 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[28]}),
		.sram(mux_tree_tapbuf_size3_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_21_sram_inv[0:1]),
		.out(chany_top_out[27]));

	mux_tree_tapbuf_size3 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[29]}),
		.sram(mux_tree_tapbuf_size3_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_22_sram_inv[0:1]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size3 mux_top_track_58 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[30]}),
		.sram(mux_tree_tapbuf_size3_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_23_sram_inv[0:1]),
		.out(chany_top_out[29]));

	mux_tree_tapbuf_size3 mux_top_track_60 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[31]}),
		.sram(mux_tree_tapbuf_size3_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_24_sram_inv[0:1]),
		.out(chany_top_out[30]));

	mux_tree_tapbuf_size3 mux_top_track_62 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[32]}),
		.sram(mux_tree_tapbuf_size3_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_25_sram_inv[0:1]),
		.out(chany_top_out[31]));

	mux_tree_tapbuf_size3 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[33]}),
		.sram(mux_tree_tapbuf_size3_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_26_sram_inv[0:1]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size3 mux_top_track_66 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[34]}),
		.sram(mux_tree_tapbuf_size3_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_27_sram_inv[0:1]),
		.out(chany_top_out[33]));

	mux_tree_tapbuf_size3 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[37]}),
		.sram(mux_tree_tapbuf_size3_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_28_sram_inv[0:1]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size3 mux_top_track_74 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[38]}),
		.sram(mux_tree_tapbuf_size3_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_29_sram_inv[0:1]),
		.out(chany_top_out[37]));

	mux_tree_tapbuf_size3 mux_top_track_76 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[39]}),
		.sram(mux_tree_tapbuf_size3_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_30_sram_inv[0:1]),
		.out(chany_top_out[38]));

	mux_tree_tapbuf_size3 mux_top_track_78 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[40]}),
		.sram(mux_tree_tapbuf_size3_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_31_sram_inv[0:1]),
		.out(chany_top_out[39]));

	mux_tree_tapbuf_size3 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[41]}),
		.sram(mux_tree_tapbuf_size3_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_32_sram_inv[0:1]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size3 mux_top_track_82 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[42]}),
		.sram(mux_tree_tapbuf_size3_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_33_sram_inv[0:1]),
		.out(chany_top_out[41]));

	mux_tree_tapbuf_size3 mux_top_track_84 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[43]}),
		.sram(mux_tree_tapbuf_size3_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_34_sram_inv[0:1]),
		.out(chany_top_out[42]));

	mux_tree_tapbuf_size3 mux_top_track_90 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[46]}),
		.sram(mux_tree_tapbuf_size3_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_35_sram_inv[0:1]),
		.out(chany_top_out[45]));

	mux_tree_tapbuf_size3 mux_top_track_92 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[47]}),
		.sram(mux_tree_tapbuf_size3_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_36_sram_inv[0:1]),
		.out(chany_top_out[46]));

	mux_tree_tapbuf_size3 mux_top_track_94 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[48]}),
		.sram(mux_tree_tapbuf_size3_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_37_sram_inv[0:1]),
		.out(chany_top_out[47]));

	mux_tree_tapbuf_size3 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[49]}),
		.sram(mux_tree_tapbuf_size3_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_38_sram_inv[0:1]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size3 mux_top_track_98 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[50]}),
		.sram(mux_tree_tapbuf_size3_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_39_sram_inv[0:1]),
		.out(chany_top_out[49]));

	mux_tree_tapbuf_size3 mux_top_track_100 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[51]}),
		.sram(mux_tree_tapbuf_size3_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_40_sram_inv[0:1]),
		.out(chany_top_out[50]));

	mux_tree_tapbuf_size3 mux_top_track_102 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[52]}),
		.sram(mux_tree_tapbuf_size3_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_41_sram_inv[0:1]),
		.out(chany_top_out[51]));

	mux_tree_tapbuf_size3 mux_top_track_108 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_size3_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_42_sram_inv[0:1]),
		.out(chany_top_out[54]));

	mux_tree_tapbuf_size3 mux_top_track_110 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_size3_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_43_sram_inv[0:1]),
		.out(chany_top_out[55]));

	mux_tree_tapbuf_size3 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_size3_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_44_sram_inv[0:1]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size3 mux_top_track_114 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[58]}),
		.sram(mux_tree_tapbuf_size3_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_45_sram_inv[0:1]),
		.out(chany_top_out[57]));

	mux_tree_tapbuf_size3 mux_top_track_116 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_size3_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_46_sram_inv[0:1]),
		.out(chany_top_out[58]));

	mux_tree_tapbuf_size3 mux_top_track_118 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_size3_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_47_sram_inv[0:1]),
		.out(chany_top_out[59]));

	mux_tree_tapbuf_size3 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_size3_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_48_sram_inv[0:1]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size3 mux_top_track_126 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_size3_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_49_sram_inv[0:1]),
		.out(chany_top_out[63]));

	mux_tree_tapbuf_size3 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_size3_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_50_sram_inv[0:1]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size3 mux_top_track_130 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[66]}),
		.sram(mux_tree_tapbuf_size3_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_51_sram_inv[0:1]),
		.out(chany_top_out[65]));

	mux_tree_tapbuf_size3 mux_top_track_132 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_size3_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_52_sram_inv[0:1]),
		.out(chany_top_out[66]));

	mux_tree_tapbuf_size3 mux_top_track_134 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_size3_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_53_sram_inv[0:1]),
		.out(chany_top_out[67]));

	mux_tree_tapbuf_size3 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_size3_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_54_sram_inv[0:1]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size3 mux_top_track_138 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[70]}),
		.sram(mux_tree_tapbuf_size3_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_55_sram_inv[0:1]),
		.out(chany_top_out[69]));

	mux_tree_tapbuf_size3 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[73]}),
		.sram(mux_tree_tapbuf_size3_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_56_sram_inv[0:1]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size3 mux_top_track_146 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[74]}),
		.sram(mux_tree_tapbuf_size3_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_57_sram_inv[0:1]),
		.out(chany_top_out[73]));

	mux_tree_tapbuf_size3 mux_top_track_148 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[75]}),
		.sram(mux_tree_tapbuf_size3_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_58_sram_inv[0:1]),
		.out(chany_top_out[74]));

	mux_tree_tapbuf_size3 mux_top_track_150 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[76]}),
		.sram(mux_tree_tapbuf_size3_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_59_sram_inv[0:1]),
		.out(chany_top_out[75]));

	mux_tree_tapbuf_size3 mux_top_track_152 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[77]}),
		.sram(mux_tree_tapbuf_size3_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_60_sram_inv[0:1]),
		.out(chany_top_out[76]));

	mux_tree_tapbuf_size3 mux_top_track_154 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[78]}),
		.sram(mux_tree_tapbuf_size3_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_61_sram_inv[0:1]),
		.out(chany_top_out[77]));

	mux_tree_tapbuf_size3 mux_top_track_156 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[79]}),
		.sram(mux_tree_tapbuf_size3_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_62_sram_inv[0:1]),
		.out(chany_top_out[78]));

	mux_tree_tapbuf_size3 mux_top_track_162 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[82]}),
		.sram(mux_tree_tapbuf_size3_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_63_sram_inv[0:1]),
		.out(chany_top_out[81]));

	mux_tree_tapbuf_size3 mux_top_track_164 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[83]}),
		.sram(mux_tree_tapbuf_size3_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_64_sram_inv[0:1]),
		.out(chany_top_out[82]));

	mux_tree_tapbuf_size3 mux_top_track_166 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[84]}),
		.sram(mux_tree_tapbuf_size3_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_65_sram_inv[0:1]),
		.out(chany_top_out[83]));

	mux_tree_tapbuf_size3 mux_top_track_168 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[85]}),
		.sram(mux_tree_tapbuf_size3_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_66_sram_inv[0:1]),
		.out(chany_top_out[84]));

	mux_tree_tapbuf_size3 mux_top_track_170 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[86]}),
		.sram(mux_tree_tapbuf_size3_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_67_sram_inv[0:1]),
		.out(chany_top_out[85]));

	mux_tree_tapbuf_size3 mux_top_track_172 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[87]}),
		.sram(mux_tree_tapbuf_size3_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_68_sram_inv[0:1]),
		.out(chany_top_out[86]));

	mux_tree_tapbuf_size3 mux_top_track_174 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[88]}),
		.sram(mux_tree_tapbuf_size3_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_69_sram_inv[0:1]),
		.out(chany_top_out[87]));

	mux_tree_tapbuf_size3 mux_top_track_180 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[91]}),
		.sram(mux_tree_tapbuf_size3_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_70_sram_inv[0:1]),
		.out(chany_top_out[90]));

	mux_tree_tapbuf_size3 mux_top_track_182 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[92]}),
		.sram(mux_tree_tapbuf_size3_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_71_sram_inv[0:1]),
		.out(chany_top_out[91]));

	mux_tree_tapbuf_size3 mux_top_track_184 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[93]}),
		.sram(mux_tree_tapbuf_size3_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_72_sram_inv[0:1]),
		.out(chany_top_out[92]));

	mux_tree_tapbuf_size3 mux_top_track_186 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[94]}),
		.sram(mux_tree_tapbuf_size3_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_73_sram_inv[0:1]),
		.out(chany_top_out[93]));

	mux_tree_tapbuf_size3 mux_top_track_188 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[95]}),
		.sram(mux_tree_tapbuf_size3_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_74_sram_inv[0:1]),
		.out(chany_top_out[94]));

	mux_tree_tapbuf_size3 mux_top_track_190 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[96]}),
		.sram(mux_tree_tapbuf_size3_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_75_sram_inv[0:1]),
		.out(chany_top_out[95]));

	mux_tree_tapbuf_size3 mux_top_track_192 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[97]}),
		.sram(mux_tree_tapbuf_size3_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_76_sram_inv[0:1]),
		.out(chany_top_out[96]));

	mux_tree_tapbuf_size3 mux_top_track_198 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[100]}),
		.sram(mux_tree_tapbuf_size3_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_77_sram_inv[0:1]),
		.out(chany_top_out[99]));

	mux_tree_tapbuf_size3 mux_top_track_200 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[101]}),
		.sram(mux_tree_tapbuf_size3_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_78_sram_inv[0:1]),
		.out(chany_top_out[100]));

	mux_tree_tapbuf_size3 mux_top_track_202 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[102]}),
		.sram(mux_tree_tapbuf_size3_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_79_sram_inv[0:1]),
		.out(chany_top_out[101]));

	mux_tree_tapbuf_size3 mux_top_track_204 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[103]}),
		.sram(mux_tree_tapbuf_size3_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_80_sram_inv[0:1]),
		.out(chany_top_out[102]));

	mux_tree_tapbuf_size3 mux_top_track_206 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[104]}),
		.sram(mux_tree_tapbuf_size3_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_81_sram_inv[0:1]),
		.out(chany_top_out[103]));

	mux_tree_tapbuf_size3 mux_top_track_208 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[105]}),
		.sram(mux_tree_tapbuf_size3_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_82_sram_inv[0:1]),
		.out(chany_top_out[104]));

	mux_tree_tapbuf_size3 mux_top_track_210 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[106]}),
		.sram(mux_tree_tapbuf_size3_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_83_sram_inv[0:1]),
		.out(chany_top_out[105]));

	mux_tree_tapbuf_size3 mux_top_track_216 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[109]}),
		.sram(mux_tree_tapbuf_size3_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_84_sram_inv[0:1]),
		.out(chany_top_out[108]));

	mux_tree_tapbuf_size3 mux_top_track_218 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[110]}),
		.sram(mux_tree_tapbuf_size3_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_85_sram_inv[0:1]),
		.out(chany_top_out[109]));

	mux_tree_tapbuf_size3 mux_top_track_220 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[111]}),
		.sram(mux_tree_tapbuf_size3_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_86_sram_inv[0:1]),
		.out(chany_top_out[110]));

	mux_tree_tapbuf_size3 mux_top_track_222 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[112]}),
		.sram(mux_tree_tapbuf_size3_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_87_sram_inv[0:1]),
		.out(chany_top_out[111]));

	mux_tree_tapbuf_size3 mux_top_track_224 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[113]}),
		.sram(mux_tree_tapbuf_size3_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_88_sram_inv[0:1]),
		.out(chany_top_out[112]));

	mux_tree_tapbuf_size3 mux_top_track_226 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[114]}),
		.sram(mux_tree_tapbuf_size3_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_89_sram_inv[0:1]),
		.out(chany_top_out[113]));

	mux_tree_tapbuf_size3 mux_top_track_228 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[115]}),
		.sram(mux_tree_tapbuf_size3_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_90_sram_inv[0:1]),
		.out(chany_top_out[114]));

	mux_tree_tapbuf_size3 mux_top_track_234 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[118]}),
		.sram(mux_tree_tapbuf_size3_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_91_sram_inv[0:1]),
		.out(chany_top_out[117]));

	mux_tree_tapbuf_size3 mux_top_track_236 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[119]}),
		.sram(mux_tree_tapbuf_size3_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_92_sram_inv[0:1]),
		.out(chany_top_out[118]));

	mux_tree_tapbuf_size3 mux_top_track_238 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[120]}),
		.sram(mux_tree_tapbuf_size3_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_93_sram_inv[0:1]),
		.out(chany_top_out[119]));

	mux_tree_tapbuf_size3 mux_top_track_240 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[121]}),
		.sram(mux_tree_tapbuf_size3_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_94_sram_inv[0:1]),
		.out(chany_top_out[120]));

	mux_tree_tapbuf_size3 mux_top_track_242 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[122]}),
		.sram(mux_tree_tapbuf_size3_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_95_sram_inv[0:1]),
		.out(chany_top_out[121]));

	mux_tree_tapbuf_size3 mux_top_track_244 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[123]}),
		.sram(mux_tree_tapbuf_size3_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_96_sram_inv[0:1]),
		.out(chany_top_out[122]));

	mux_tree_tapbuf_size3 mux_top_track_246 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[124]}),
		.sram(mux_tree_tapbuf_size3_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_97_sram_inv[0:1]),
		.out(chany_top_out[123]));

	mux_tree_tapbuf_size3 mux_top_track_252 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[127]}),
		.sram(mux_tree_tapbuf_size3_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_98_sram_inv[0:1]),
		.out(chany_top_out[126]));

	mux_tree_tapbuf_size3 mux_top_track_254 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[128]}),
		.sram(mux_tree_tapbuf_size3_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_99_sram_inv[0:1]),
		.out(chany_top_out[127]));

	mux_tree_tapbuf_size3 mux_top_track_256 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[129]}),
		.sram(mux_tree_tapbuf_size3_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_100_sram_inv[0:1]),
		.out(chany_top_out[128]));

	mux_tree_tapbuf_size3 mux_top_track_258 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[130]}),
		.sram(mux_tree_tapbuf_size3_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_101_sram_inv[0:1]),
		.out(chany_top_out[129]));

	mux_tree_tapbuf_size3 mux_top_track_260 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[131]}),
		.sram(mux_tree_tapbuf_size3_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_102_sram_inv[0:1]),
		.out(chany_top_out[130]));

	mux_tree_tapbuf_size3 mux_top_track_262 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[132]}),
		.sram(mux_tree_tapbuf_size3_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_103_sram_inv[0:1]),
		.out(chany_top_out[131]));

	mux_tree_tapbuf_size3 mux_top_track_264 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[133]}),
		.sram(mux_tree_tapbuf_size3_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_104_sram_inv[0:1]),
		.out(chany_top_out[132]));

	mux_tree_tapbuf_size3 mux_top_track_270 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[136]}),
		.sram(mux_tree_tapbuf_size3_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_105_sram_inv[0:1]),
		.out(chany_top_out[135]));

	mux_tree_tapbuf_size3 mux_top_track_272 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[137]}),
		.sram(mux_tree_tapbuf_size3_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_106_sram_inv[0:1]),
		.out(chany_top_out[136]));

	mux_tree_tapbuf_size3 mux_top_track_274 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[138]}),
		.sram(mux_tree_tapbuf_size3_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_107_sram_inv[0:1]),
		.out(chany_top_out[137]));

	mux_tree_tapbuf_size3 mux_top_track_276 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[139]}),
		.sram(mux_tree_tapbuf_size3_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_108_sram_inv[0:1]),
		.out(chany_top_out[138]));

	mux_tree_tapbuf_size3 mux_top_track_278 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[140]}),
		.sram(mux_tree_tapbuf_size3_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_109_sram_inv[0:1]),
		.out(chany_top_out[139]));

	mux_tree_tapbuf_size3 mux_top_track_280 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[141]}),
		.sram(mux_tree_tapbuf_size3_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_110_sram_inv[0:1]),
		.out(chany_top_out[140]));

	mux_tree_tapbuf_size3 mux_top_track_282 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[142]}),
		.sram(mux_tree_tapbuf_size3_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_111_sram_inv[0:1]),
		.out(chany_top_out[141]));

	mux_tree_tapbuf_size3 mux_top_track_288 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[145]}),
		.sram(mux_tree_tapbuf_size3_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_112_sram_inv[0:1]),
		.out(chany_top_out[144]));

	mux_tree_tapbuf_size3 mux_top_track_290 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[146]}),
		.sram(mux_tree_tapbuf_size3_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_113_sram_inv[0:1]),
		.out(chany_top_out[145]));

	mux_tree_tapbuf_size3 mux_top_track_292 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[147]}),
		.sram(mux_tree_tapbuf_size3_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_114_sram_inv[0:1]),
		.out(chany_top_out[146]));

	mux_tree_tapbuf_size3 mux_top_track_294 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[148]}),
		.sram(mux_tree_tapbuf_size3_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_115_sram_inv[0:1]),
		.out(chany_top_out[147]));

	mux_tree_tapbuf_size3 mux_top_track_296 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[149]}),
		.sram(mux_tree_tapbuf_size3_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_116_sram_inv[0:1]),
		.out(chany_top_out[148]));

	mux_tree_tapbuf_size3 mux_top_track_298 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[150]}),
		.sram(mux_tree_tapbuf_size3_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_117_sram_inv[0:1]),
		.out(chany_top_out[149]));

	mux_tree_tapbuf_size3 mux_top_track_300 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[151]}),
		.sram(mux_tree_tapbuf_size3_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_118_sram_inv[0:1]),
		.out(chany_top_out[150]));

	mux_tree_tapbuf_size3 mux_top_track_306 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[154]}),
		.sram(mux_tree_tapbuf_size3_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_119_sram_inv[0:1]),
		.out(chany_top_out[153]));

	mux_tree_tapbuf_size3 mux_top_track_308 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[155]}),
		.sram(mux_tree_tapbuf_size3_120_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_120_sram_inv[0:1]),
		.out(chany_top_out[154]));

	mux_tree_tapbuf_size3 mux_top_track_310 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[156]}),
		.sram(mux_tree_tapbuf_size3_121_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_121_sram_inv[0:1]),
		.out(chany_top_out[155]));

	mux_tree_tapbuf_size3 mux_top_track_312 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[157]}),
		.sram(mux_tree_tapbuf_size3_122_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_122_sram_inv[0:1]),
		.out(chany_top_out[156]));

	mux_tree_tapbuf_size3 mux_top_track_314 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[158]}),
		.sram(mux_tree_tapbuf_size3_123_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_123_sram_inv[0:1]),
		.out(chany_top_out[157]));

	mux_tree_tapbuf_size3 mux_top_track_316 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[159]}),
		.sram(mux_tree_tapbuf_size3_124_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_124_sram_inv[0:1]),
		.out(chany_top_out[158]));

	mux_tree_tapbuf_size3 mux_top_track_318 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[160]}),
		.sram(mux_tree_tapbuf_size3_125_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_125_sram_inv[0:1]),
		.out(chany_top_out[159]));

	mux_tree_tapbuf_size3 mux_top_track_324 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[163]}),
		.sram(mux_tree_tapbuf_size3_126_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_126_sram_inv[0:1]),
		.out(chany_top_out[162]));

	mux_tree_tapbuf_size3 mux_top_track_326 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[164]}),
		.sram(mux_tree_tapbuf_size3_127_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_127_sram_inv[0:1]),
		.out(chany_top_out[163]));

	mux_tree_tapbuf_size3 mux_top_track_328 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[165]}),
		.sram(mux_tree_tapbuf_size3_128_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_128_sram_inv[0:1]),
		.out(chany_top_out[164]));

	mux_tree_tapbuf_size3 mux_top_track_330 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[166]}),
		.sram(mux_tree_tapbuf_size3_129_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_129_sram_inv[0:1]),
		.out(chany_top_out[165]));

	mux_tree_tapbuf_size3 mux_top_track_332 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[167]}),
		.sram(mux_tree_tapbuf_size3_130_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_130_sram_inv[0:1]),
		.out(chany_top_out[166]));

	mux_tree_tapbuf_size3 mux_top_track_334 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[168]}),
		.sram(mux_tree_tapbuf_size3_131_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_131_sram_inv[0:1]),
		.out(chany_top_out[167]));

	mux_tree_tapbuf_size3 mux_top_track_336 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[169]}),
		.sram(mux_tree_tapbuf_size3_132_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_132_sram_inv[0:1]),
		.out(chany_top_out[168]));

	mux_tree_tapbuf_size3 mux_top_track_342 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[172]}),
		.sram(mux_tree_tapbuf_size3_133_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_133_sram_inv[0:1]),
		.out(chany_top_out[171]));

	mux_tree_tapbuf_size3 mux_top_track_344 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[173]}),
		.sram(mux_tree_tapbuf_size3_134_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_134_sram_inv[0:1]),
		.out(chany_top_out[172]));

	mux_tree_tapbuf_size3 mux_top_track_346 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[174]}),
		.sram(mux_tree_tapbuf_size3_135_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_135_sram_inv[0:1]),
		.out(chany_top_out[173]));

	mux_tree_tapbuf_size3 mux_top_track_348 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[175]}),
		.sram(mux_tree_tapbuf_size3_136_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_136_sram_inv[0:1]),
		.out(chany_top_out[174]));

	mux_tree_tapbuf_size3 mux_top_track_350 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[176]}),
		.sram(mux_tree_tapbuf_size3_137_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_137_sram_inv[0:1]),
		.out(chany_top_out[175]));

	mux_tree_tapbuf_size3 mux_top_track_352 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[177]}),
		.sram(mux_tree_tapbuf_size3_138_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_138_sram_inv[0:1]),
		.out(chany_top_out[176]));

	mux_tree_tapbuf_size3 mux_top_track_354 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[178]}),
		.sram(mux_tree_tapbuf_size3_139_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_139_sram_inv[0:1]),
		.out(chany_top_out[177]));

	mux_tree_tapbuf_size3 mux_top_track_360 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[181]}),
		.sram(mux_tree_tapbuf_size3_140_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_140_sram_inv[0:1]),
		.out(chany_top_out[180]));

	mux_tree_tapbuf_size3 mux_top_track_362 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[182]}),
		.sram(mux_tree_tapbuf_size3_141_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_141_sram_inv[0:1]),
		.out(chany_top_out[181]));

	mux_tree_tapbuf_size3 mux_top_track_364 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[183]}),
		.sram(mux_tree_tapbuf_size3_142_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_142_sram_inv[0:1]),
		.out(chany_top_out[182]));

	mux_tree_tapbuf_size3 mux_top_track_366 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[184]}),
		.sram(mux_tree_tapbuf_size3_143_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_143_sram_inv[0:1]),
		.out(chany_top_out[183]));

	mux_tree_tapbuf_size3 mux_top_track_368 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[185]}),
		.sram(mux_tree_tapbuf_size3_144_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_144_sram_inv[0:1]),
		.out(chany_top_out[184]));

	mux_tree_tapbuf_size3 mux_top_track_370 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[186]}),
		.sram(mux_tree_tapbuf_size3_145_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_145_sram_inv[0:1]),
		.out(chany_top_out[185]));

	mux_tree_tapbuf_size3 mux_top_track_372 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[187]}),
		.sram(mux_tree_tapbuf_size3_146_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_146_sram_inv[0:1]),
		.out(chany_top_out[186]));

	mux_tree_tapbuf_size3 mux_top_track_378 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[190]}),
		.sram(mux_tree_tapbuf_size3_147_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_147_sram_inv[0:1]),
		.out(chany_top_out[189]));

	mux_tree_tapbuf_size3 mux_top_track_380 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[191]}),
		.sram(mux_tree_tapbuf_size3_148_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_148_sram_inv[0:1]),
		.out(chany_top_out[190]));

	mux_tree_tapbuf_size3 mux_top_track_382 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[192]}),
		.sram(mux_tree_tapbuf_size3_149_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_149_sram_inv[0:1]),
		.out(chany_top_out[191]));

	mux_tree_tapbuf_size3 mux_top_track_384 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[193]}),
		.sram(mux_tree_tapbuf_size3_150_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_150_sram_inv[0:1]),
		.out(chany_top_out[192]));

	mux_tree_tapbuf_size3 mux_top_track_386 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[194]}),
		.sram(mux_tree_tapbuf_size3_151_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_151_sram_inv[0:1]),
		.out(chany_top_out[193]));

	mux_tree_tapbuf_size3 mux_top_track_388 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[195]}),
		.sram(mux_tree_tapbuf_size3_152_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_152_sram_inv[0:1]),
		.out(chany_top_out[194]));

	mux_tree_tapbuf_size3 mux_top_track_390 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[196]}),
		.sram(mux_tree_tapbuf_size3_153_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_153_sram_inv[0:1]),
		.out(chany_top_out[195]));

	mux_tree_tapbuf_size3 mux_top_track_396 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[199]}),
		.sram(mux_tree_tapbuf_size3_154_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_154_sram_inv[0:1]),
		.out(chany_top_out[198]));

	mux_tree_tapbuf_size3 mux_top_track_398 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[200]}),
		.sram(mux_tree_tapbuf_size3_155_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_155_sram_inv[0:1]),
		.out(chany_top_out[199]));

	mux_tree_tapbuf_size3 mux_top_track_400 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[201]}),
		.sram(mux_tree_tapbuf_size3_156_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_156_sram_inv[0:1]),
		.out(chany_top_out[200]));

	mux_tree_tapbuf_size3 mux_top_track_402 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[202]}),
		.sram(mux_tree_tapbuf_size3_157_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_157_sram_inv[0:1]),
		.out(chany_top_out[201]));

	mux_tree_tapbuf_size3 mux_top_track_404 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[203]}),
		.sram(mux_tree_tapbuf_size3_158_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_158_sram_inv[0:1]),
		.out(chany_top_out[202]));

	mux_tree_tapbuf_size3 mux_top_track_406 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[204]}),
		.sram(mux_tree_tapbuf_size3_159_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_159_sram_inv[0:1]),
		.out(chany_top_out[203]));

	mux_tree_tapbuf_size3 mux_top_track_408 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[205]}),
		.sram(mux_tree_tapbuf_size3_160_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_160_sram_inv[0:1]),
		.out(chany_top_out[204]));

	mux_tree_tapbuf_size3 mux_top_track_414 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[208]}),
		.sram(mux_tree_tapbuf_size3_161_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_161_sram_inv[0:1]),
		.out(chany_top_out[207]));

	mux_tree_tapbuf_size3 mux_top_track_416 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[209]}),
		.sram(mux_tree_tapbuf_size3_162_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_162_sram_inv[0:1]),
		.out(chany_top_out[208]));

	mux_tree_tapbuf_size3 mux_top_track_418 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[210]}),
		.sram(mux_tree_tapbuf_size3_163_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_163_sram_inv[0:1]),
		.out(chany_top_out[209]));

	mux_tree_tapbuf_size3 mux_top_track_420 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[211]}),
		.sram(mux_tree_tapbuf_size3_164_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_164_sram_inv[0:1]),
		.out(chany_top_out[210]));

	mux_tree_tapbuf_size3 mux_top_track_422 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[212]}),
		.sram(mux_tree_tapbuf_size3_165_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_165_sram_inv[0:1]),
		.out(chany_top_out[211]));

	mux_tree_tapbuf_size3 mux_top_track_424 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[213]}),
		.sram(mux_tree_tapbuf_size3_166_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_166_sram_inv[0:1]),
		.out(chany_top_out[212]));

	mux_tree_tapbuf_size3 mux_top_track_426 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[214]}),
		.sram(mux_tree_tapbuf_size3_167_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_167_sram_inv[0:1]),
		.out(chany_top_out[213]));

	mux_tree_tapbuf_size3 mux_top_track_432 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[217]}),
		.sram(mux_tree_tapbuf_size3_168_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_168_sram_inv[0:1]),
		.out(chany_top_out[216]));

	mux_tree_tapbuf_size3 mux_top_track_434 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[218]}),
		.sram(mux_tree_tapbuf_size3_169_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_169_sram_inv[0:1]),
		.out(chany_top_out[217]));

	mux_tree_tapbuf_size3 mux_top_track_436 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[219]}),
		.sram(mux_tree_tapbuf_size3_170_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_170_sram_inv[0:1]),
		.out(chany_top_out[218]));

	mux_tree_tapbuf_size3 mux_top_track_438 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[220]}),
		.sram(mux_tree_tapbuf_size3_171_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_171_sram_inv[0:1]),
		.out(chany_top_out[219]));

	mux_tree_tapbuf_size3 mux_top_track_440 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[221]}),
		.sram(mux_tree_tapbuf_size3_172_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_172_sram_inv[0:1]),
		.out(chany_top_out[220]));

	mux_tree_tapbuf_size3 mux_top_track_442 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[222]}),
		.sram(mux_tree_tapbuf_size3_173_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_173_sram_inv[0:1]),
		.out(chany_top_out[221]));

	mux_tree_tapbuf_size3 mux_top_track_444 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[223]}),
		.sram(mux_tree_tapbuf_size3_174_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_174_sram_inv[0:1]),
		.out(chany_top_out[222]));

	mux_tree_tapbuf_size3 mux_top_track_450 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[226]}),
		.sram(mux_tree_tapbuf_size3_175_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_175_sram_inv[0:1]),
		.out(chany_top_out[225]));

	mux_tree_tapbuf_size3 mux_top_track_452 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[227]}),
		.sram(mux_tree_tapbuf_size3_176_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_176_sram_inv[0:1]),
		.out(chany_top_out[226]));

	mux_tree_tapbuf_size3 mux_top_track_454 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[228]}),
		.sram(mux_tree_tapbuf_size3_177_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_177_sram_inv[0:1]),
		.out(chany_top_out[227]));

	mux_tree_tapbuf_size3 mux_top_track_456 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[229]}),
		.sram(mux_tree_tapbuf_size3_178_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_178_sram_inv[0:1]),
		.out(chany_top_out[228]));

	mux_tree_tapbuf_size3 mux_top_track_458 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[230]}),
		.sram(mux_tree_tapbuf_size3_179_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_179_sram_inv[0:1]),
		.out(chany_top_out[229]));

	mux_tree_tapbuf_size3 mux_top_track_460 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[231]}),
		.sram(mux_tree_tapbuf_size3_180_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_180_sram_inv[0:1]),
		.out(chany_top_out[230]));

	mux_tree_tapbuf_size3 mux_top_track_462 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[232]}),
		.sram(mux_tree_tapbuf_size3_181_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_181_sram_inv[0:1]),
		.out(chany_top_out[231]));

	mux_tree_tapbuf_size3 mux_top_track_468 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[235]}),
		.sram(mux_tree_tapbuf_size3_182_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_182_sram_inv[0:1]),
		.out(chany_top_out[234]));

	mux_tree_tapbuf_size3 mux_top_track_470 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[236]}),
		.sram(mux_tree_tapbuf_size3_183_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_183_sram_inv[0:1]),
		.out(chany_top_out[235]));

	mux_tree_tapbuf_size3 mux_top_track_472 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[237]}),
		.sram(mux_tree_tapbuf_size3_184_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_184_sram_inv[0:1]),
		.out(chany_top_out[236]));

	mux_tree_tapbuf_size3 mux_top_track_474 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[238]}),
		.sram(mux_tree_tapbuf_size3_185_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_185_sram_inv[0:1]),
		.out(chany_top_out[237]));

	mux_tree_tapbuf_size3 mux_top_track_476 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[239]}),
		.sram(mux_tree_tapbuf_size3_186_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_186_sram_inv[0:1]),
		.out(chany_top_out[238]));

	mux_tree_tapbuf_size3 mux_top_track_478 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[240]}),
		.sram(mux_tree_tapbuf_size3_187_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_187_sram_inv[0:1]),
		.out(chany_top_out[239]));

	mux_tree_tapbuf_size3 mux_top_track_480 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[241]}),
		.sram(mux_tree_tapbuf_size3_188_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_188_sram_inv[0:1]),
		.out(chany_top_out[240]));

	mux_tree_tapbuf_size3 mux_top_track_486 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[244]}),
		.sram(mux_tree_tapbuf_size3_189_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_189_sram_inv[0:1]),
		.out(chany_top_out[243]));

	mux_tree_tapbuf_size3 mux_top_track_488 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[245]}),
		.sram(mux_tree_tapbuf_size3_190_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_190_sram_inv[0:1]),
		.out(chany_top_out[244]));

	mux_tree_tapbuf_size3 mux_top_track_490 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[246]}),
		.sram(mux_tree_tapbuf_size3_191_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_191_sram_inv[0:1]),
		.out(chany_top_out[245]));

	mux_tree_tapbuf_size3 mux_top_track_492 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[247]}),
		.sram(mux_tree_tapbuf_size3_192_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_192_sram_inv[0:1]),
		.out(chany_top_out[246]));

	mux_tree_tapbuf_size3 mux_top_track_494 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[248]}),
		.sram(mux_tree_tapbuf_size3_193_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_193_sram_inv[0:1]),
		.out(chany_top_out[247]));

	mux_tree_tapbuf_size3 mux_top_track_496 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[249]}),
		.sram(mux_tree_tapbuf_size3_194_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_194_sram_inv[0:1]),
		.out(chany_top_out[248]));

	mux_tree_tapbuf_size3 mux_top_track_498 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[250]}),
		.sram(mux_tree_tapbuf_size3_195_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_195_sram_inv[0:1]),
		.out(chany_top_out[249]));

	mux_tree_tapbuf_size3 mux_top_track_504 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[253]}),
		.sram(mux_tree_tapbuf_size3_196_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_196_sram_inv[0:1]),
		.out(chany_top_out[252]));

	mux_tree_tapbuf_size3 mux_top_track_506 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[254]}),
		.sram(mux_tree_tapbuf_size3_197_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_197_sram_inv[0:1]),
		.out(chany_top_out[253]));

	mux_tree_tapbuf_size3 mux_top_track_508 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[255]}),
		.sram(mux_tree_tapbuf_size3_198_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_198_sram_inv[0:1]),
		.out(chany_top_out[254]));

	mux_tree_tapbuf_size3 mux_top_track_510 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[256]}),
		.sram(mux_tree_tapbuf_size3_199_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_199_sram_inv[0:1]),
		.out(chany_top_out[255]));

	mux_tree_tapbuf_size3 mux_top_track_512 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[257]}),
		.sram(mux_tree_tapbuf_size3_200_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_200_sram_inv[0:1]),
		.out(chany_top_out[256]));

	mux_tree_tapbuf_size3 mux_top_track_514 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[258]}),
		.sram(mux_tree_tapbuf_size3_201_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_201_sram_inv[0:1]),
		.out(chany_top_out[257]));

	mux_tree_tapbuf_size3 mux_top_track_516 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[259]}),
		.sram(mux_tree_tapbuf_size3_202_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_202_sram_inv[0:1]),
		.out(chany_top_out[258]));

	mux_tree_tapbuf_size3 mux_top_track_522 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[262]}),
		.sram(mux_tree_tapbuf_size3_203_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_203_sram_inv[0:1]),
		.out(chany_top_out[261]));

	mux_tree_tapbuf_size3 mux_top_track_524 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[263]}),
		.sram(mux_tree_tapbuf_size3_204_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_204_sram_inv[0:1]),
		.out(chany_top_out[262]));

	mux_tree_tapbuf_size3 mux_top_track_526 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[264]}),
		.sram(mux_tree_tapbuf_size3_205_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_205_sram_inv[0:1]),
		.out(chany_top_out[263]));

	mux_tree_tapbuf_size3 mux_top_track_528 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[265]}),
		.sram(mux_tree_tapbuf_size3_206_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_206_sram_inv[0:1]),
		.out(chany_top_out[264]));

	mux_tree_tapbuf_size3 mux_top_track_530 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[266]}),
		.sram(mux_tree_tapbuf_size3_207_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_207_sram_inv[0:1]),
		.out(chany_top_out[265]));

	mux_tree_tapbuf_size3 mux_top_track_532 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[267]}),
		.sram(mux_tree_tapbuf_size3_208_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_208_sram_inv[0:1]),
		.out(chany_top_out[266]));

	mux_tree_tapbuf_size3 mux_top_track_534 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[268]}),
		.sram(mux_tree_tapbuf_size3_209_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_209_sram_inv[0:1]),
		.out(chany_top_out[267]));

	mux_tree_tapbuf_size3 mux_top_track_540 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[271]}),
		.sram(mux_tree_tapbuf_size3_210_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_210_sram_inv[0:1]),
		.out(chany_top_out[270]));

	mux_tree_tapbuf_size3 mux_top_track_542 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[272]}),
		.sram(mux_tree_tapbuf_size3_211_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_211_sram_inv[0:1]),
		.out(chany_top_out[271]));

	mux_tree_tapbuf_size3 mux_top_track_544 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[273]}),
		.sram(mux_tree_tapbuf_size3_212_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_212_sram_inv[0:1]),
		.out(chany_top_out[272]));

	mux_tree_tapbuf_size3 mux_top_track_546 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[274]}),
		.sram(mux_tree_tapbuf_size3_213_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_213_sram_inv[0:1]),
		.out(chany_top_out[273]));

	mux_tree_tapbuf_size3 mux_top_track_548 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[275]}),
		.sram(mux_tree_tapbuf_size3_214_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_214_sram_inv[0:1]),
		.out(chany_top_out[274]));

	mux_tree_tapbuf_size3 mux_top_track_550 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[276]}),
		.sram(mux_tree_tapbuf_size3_215_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_215_sram_inv[0:1]),
		.out(chany_top_out[275]));

	mux_tree_tapbuf_size3 mux_top_track_552 (
		.in({top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[277]}),
		.sram(mux_tree_tapbuf_size3_216_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_216_sram_inv[0:1]),
		.out(chany_top_out[276]));

	mux_tree_tapbuf_size3 mux_top_track_558 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_, chanx_right_in[280]}),
		.sram(mux_tree_tapbuf_size3_217_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_217_sram_inv[0:1]),
		.out(chany_top_out[279]));

	mux_tree_tapbuf_size3 mux_top_track_560 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_, chanx_right_in[281]}),
		.sram(mux_tree_tapbuf_size3_218_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_218_sram_inv[0:1]),
		.out(chany_top_out[280]));

	mux_tree_tapbuf_size3 mux_top_track_562 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_, chanx_right_in[282]}),
		.sram(mux_tree_tapbuf_size3_219_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_219_sram_inv[0:1]),
		.out(chany_top_out[281]));

	mux_tree_tapbuf_size3 mux_top_track_564 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_, chanx_right_in[283]}),
		.sram(mux_tree_tapbuf_size3_220_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_220_sram_inv[0:1]),
		.out(chany_top_out[282]));

	mux_tree_tapbuf_size3 mux_top_track_566 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_, chanx_right_in[284]}),
		.sram(mux_tree_tapbuf_size3_221_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_221_sram_inv[0:1]),
		.out(chany_top_out[283]));

	mux_tree_tapbuf_size3 mux_top_track_568 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_, chanx_right_in[0]}),
		.sram(mux_tree_tapbuf_size3_222_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_222_sram_inv[0:1]),
		.out(chany_top_out[284]));

	mux_tree_tapbuf_size3 mux_right_track_2 (
		.in({chany_top_in[0], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_223_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_223_sram_inv[0:1]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size3 mux_right_track_4 (
		.in({chany_top_in[1], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_224_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_224_sram_inv[0:1]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size3 mux_right_track_6 (
		.in({chany_top_in[2], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_225_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_225_sram_inv[0:1]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size3 mux_right_track_8 (
		.in({chany_top_in[3], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_226_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_226_sram_inv[0:1]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size3 mux_right_track_10 (
		.in({chany_top_in[4], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_227_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_227_sram_inv[0:1]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size3 mux_right_track_12 (
		.in({chany_top_in[5], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_228_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_228_sram_inv[0:1]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size3 mux_right_track_14 (
		.in({chany_top_in[6], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_229_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_229_sram_inv[0:1]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size3 mux_right_track_16 (
		.in({chany_top_in[7], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_230_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_230_sram_inv[0:1]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size3 mux_right_track_20 (
		.in({chany_top_in[9], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_231_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_231_sram_inv[0:1]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size3 mux_right_track_22 (
		.in({chany_top_in[10], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_232_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_232_sram_inv[0:1]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size3 mux_right_track_24 (
		.in({chany_top_in[11], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_233_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_233_sram_inv[0:1]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size3 mux_right_track_26 (
		.in({chany_top_in[12], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_234_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_234_sram_inv[0:1]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size3 mux_right_track_28 (
		.in({chany_top_in[13], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_235_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_235_sram_inv[0:1]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size3 mux_right_track_30 (
		.in({chany_top_in[14], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_236_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_236_sram_inv[0:1]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size3 mux_right_track_36 (
		.in({chany_top_in[17], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_237_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_237_sram_inv[0:1]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size3 mux_right_track_38 (
		.in({chany_top_in[18], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_238_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_238_sram_inv[0:1]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size3 mux_right_track_40 (
		.in({chany_top_in[19], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_239_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_239_sram_inv[0:1]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size3 mux_right_track_42 (
		.in({chany_top_in[20], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_240_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_240_sram_inv[0:1]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size3 mux_right_track_44 (
		.in({chany_top_in[21], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_241_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_241_sram_inv[0:1]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size3 mux_right_track_46 (
		.in({chany_top_in[22], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_242_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_242_sram_inv[0:1]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size3 mux_right_track_48 (
		.in({chany_top_in[23], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_243_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_243_sram_inv[0:1]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size3 mux_right_track_54 (
		.in({chany_top_in[26], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_244_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_244_sram_inv[0:1]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size3 mux_right_track_56 (
		.in({chany_top_in[27], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_245_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_245_sram_inv[0:1]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size3 mux_right_track_58 (
		.in({chany_top_in[28], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_246_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_246_sram_inv[0:1]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size3 mux_right_track_60 (
		.in({chany_top_in[29], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_247_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_247_sram_inv[0:1]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size3 mux_right_track_62 (
		.in({chany_top_in[30], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_248_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_248_sram_inv[0:1]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size3 mux_right_track_64 (
		.in({chany_top_in[31], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_249_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_249_sram_inv[0:1]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size3 mux_right_track_66 (
		.in({chany_top_in[32], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_250_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_250_sram_inv[0:1]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size3 mux_right_track_72 (
		.in({chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_251_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_251_sram_inv[0:1]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size3 mux_right_track_74 (
		.in({chany_top_in[36], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_252_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_252_sram_inv[0:1]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size3 mux_right_track_76 (
		.in({chany_top_in[37], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_253_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_253_sram_inv[0:1]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size3 mux_right_track_78 (
		.in({chany_top_in[38], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_254_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_254_sram_inv[0:1]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size3 mux_right_track_80 (
		.in({chany_top_in[39], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_255_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_255_sram_inv[0:1]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size3 mux_right_track_82 (
		.in({chany_top_in[40], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_256_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_256_sram_inv[0:1]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size3 mux_right_track_84 (
		.in({chany_top_in[41], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_257_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_257_sram_inv[0:1]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size3 mux_right_track_90 (
		.in({chany_top_in[44], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_258_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_258_sram_inv[0:1]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size3 mux_right_track_92 (
		.in({chany_top_in[45], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_259_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_259_sram_inv[0:1]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size3 mux_right_track_94 (
		.in({chany_top_in[46], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_260_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_260_sram_inv[0:1]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size3 mux_right_track_96 (
		.in({chany_top_in[47], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_261_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_261_sram_inv[0:1]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size3 mux_right_track_98 (
		.in({chany_top_in[48], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_262_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_262_sram_inv[0:1]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size3 mux_right_track_100 (
		.in({chany_top_in[49], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_263_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_263_sram_inv[0:1]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size3 mux_right_track_102 (
		.in({chany_top_in[50], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_264_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_264_sram_inv[0:1]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size3 mux_right_track_108 (
		.in({chany_top_in[53], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_265_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_265_sram_inv[0:1]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size3 mux_right_track_110 (
		.in({chany_top_in[54], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_266_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_266_sram_inv[0:1]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size3 mux_right_track_112 (
		.in({chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_267_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_267_sram_inv[0:1]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size3 mux_right_track_114 (
		.in({chany_top_in[56], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_268_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_268_sram_inv[0:1]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size3 mux_right_track_116 (
		.in({chany_top_in[57], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_269_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_269_sram_inv[0:1]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size3 mux_right_track_118 (
		.in({chany_top_in[58], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_270_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_270_sram_inv[0:1]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size3 mux_right_track_120 (
		.in({chany_top_in[59], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_271_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_271_sram_inv[0:1]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size3 mux_right_track_126 (
		.in({chany_top_in[62], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_272_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_272_sram_inv[0:1]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size3 mux_right_track_128 (
		.in({chany_top_in[63], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_273_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_273_sram_inv[0:1]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size3 mux_right_track_130 (
		.in({chany_top_in[64], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_274_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_274_sram_inv[0:1]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size3 mux_right_track_132 (
		.in({chany_top_in[65], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_275_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_275_sram_inv[0:1]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size3 mux_right_track_134 (
		.in({chany_top_in[66], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_276_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_276_sram_inv[0:1]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size3 mux_right_track_136 (
		.in({chany_top_in[67], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_277_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_277_sram_inv[0:1]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size3 mux_right_track_138 (
		.in({chany_top_in[68], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_278_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_278_sram_inv[0:1]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size3 mux_right_track_144 (
		.in({chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_279_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_279_sram_inv[0:1]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size3 mux_right_track_146 (
		.in({chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_280_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_280_sram_inv[0:1]),
		.out(chanx_right_out[73]));

	mux_tree_tapbuf_size3 mux_right_track_148 (
		.in({chany_top_in[73], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_281_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_281_sram_inv[0:1]),
		.out(chanx_right_out[74]));

	mux_tree_tapbuf_size3 mux_right_track_150 (
		.in({chany_top_in[74], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_282_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_282_sram_inv[0:1]),
		.out(chanx_right_out[75]));

	mux_tree_tapbuf_size3 mux_right_track_152 (
		.in({chany_top_in[75], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_283_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_283_sram_inv[0:1]),
		.out(chanx_right_out[76]));

	mux_tree_tapbuf_size3 mux_right_track_154 (
		.in({chany_top_in[76], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_284_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_284_sram_inv[0:1]),
		.out(chanx_right_out[77]));

	mux_tree_tapbuf_size3 mux_right_track_156 (
		.in({chany_top_in[77], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_285_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_285_sram_inv[0:1]),
		.out(chanx_right_out[78]));

	mux_tree_tapbuf_size3 mux_right_track_162 (
		.in({chany_top_in[80], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_286_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_286_sram_inv[0:1]),
		.out(chanx_right_out[81]));

	mux_tree_tapbuf_size3 mux_right_track_164 (
		.in({chany_top_in[81], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_287_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_287_sram_inv[0:1]),
		.out(chanx_right_out[82]));

	mux_tree_tapbuf_size3 mux_right_track_166 (
		.in({chany_top_in[82], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_288_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_288_sram_inv[0:1]),
		.out(chanx_right_out[83]));

	mux_tree_tapbuf_size3 mux_right_track_168 (
		.in({chany_top_in[83], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_289_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_289_sram_inv[0:1]),
		.out(chanx_right_out[84]));

	mux_tree_tapbuf_size3 mux_right_track_170 (
		.in({chany_top_in[84], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_290_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_290_sram_inv[0:1]),
		.out(chanx_right_out[85]));

	mux_tree_tapbuf_size3 mux_right_track_172 (
		.in({chany_top_in[85], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_291_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_291_sram_inv[0:1]),
		.out(chanx_right_out[86]));

	mux_tree_tapbuf_size3 mux_right_track_174 (
		.in({chany_top_in[86], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_292_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_292_sram_inv[0:1]),
		.out(chanx_right_out[87]));

	mux_tree_tapbuf_size3 mux_right_track_180 (
		.in({chany_top_in[89], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_293_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_293_sram_inv[0:1]),
		.out(chanx_right_out[90]));

	mux_tree_tapbuf_size3 mux_right_track_182 (
		.in({chany_top_in[90], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_294_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_294_sram_inv[0:1]),
		.out(chanx_right_out[91]));

	mux_tree_tapbuf_size3 mux_right_track_184 (
		.in({chany_top_in[91], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_295_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_295_sram_inv[0:1]),
		.out(chanx_right_out[92]));

	mux_tree_tapbuf_size3 mux_right_track_186 (
		.in({chany_top_in[92], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_296_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_296_sram_inv[0:1]),
		.out(chanx_right_out[93]));

	mux_tree_tapbuf_size3 mux_right_track_188 (
		.in({chany_top_in[93], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_297_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_297_sram_inv[0:1]),
		.out(chanx_right_out[94]));

	mux_tree_tapbuf_size3 mux_right_track_190 (
		.in({chany_top_in[94], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_298_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_298_sram_inv[0:1]),
		.out(chanx_right_out[95]));

	mux_tree_tapbuf_size3 mux_right_track_192 (
		.in({chany_top_in[95], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_299_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_299_sram_inv[0:1]),
		.out(chanx_right_out[96]));

	mux_tree_tapbuf_size3 mux_right_track_198 (
		.in({chany_top_in[98], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_300_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_300_sram_inv[0:1]),
		.out(chanx_right_out[99]));

	mux_tree_tapbuf_size3 mux_right_track_200 (
		.in({chany_top_in[99], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_301_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_301_sram_inv[0:1]),
		.out(chanx_right_out[100]));

	mux_tree_tapbuf_size3 mux_right_track_202 (
		.in({chany_top_in[100], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_302_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_302_sram_inv[0:1]),
		.out(chanx_right_out[101]));

	mux_tree_tapbuf_size3 mux_right_track_204 (
		.in({chany_top_in[101], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_303_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_303_sram_inv[0:1]),
		.out(chanx_right_out[102]));

	mux_tree_tapbuf_size3 mux_right_track_206 (
		.in({chany_top_in[102], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_304_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_304_sram_inv[0:1]),
		.out(chanx_right_out[103]));

	mux_tree_tapbuf_size3 mux_right_track_208 (
		.in({chany_top_in[103], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_305_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_305_sram_inv[0:1]),
		.out(chanx_right_out[104]));

	mux_tree_tapbuf_size3 mux_right_track_210 (
		.in({chany_top_in[104], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_306_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_306_sram_inv[0:1]),
		.out(chanx_right_out[105]));

	mux_tree_tapbuf_size3 mux_right_track_216 (
		.in({chany_top_in[107], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_307_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_307_sram_inv[0:1]),
		.out(chanx_right_out[108]));

	mux_tree_tapbuf_size3 mux_right_track_218 (
		.in({chany_top_in[108], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_308_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_308_sram_inv[0:1]),
		.out(chanx_right_out[109]));

	mux_tree_tapbuf_size3 mux_right_track_220 (
		.in({chany_top_in[109], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_309_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_309_sram_inv[0:1]),
		.out(chanx_right_out[110]));

	mux_tree_tapbuf_size3 mux_right_track_222 (
		.in({chany_top_in[110], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_310_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_310_sram_inv[0:1]),
		.out(chanx_right_out[111]));

	mux_tree_tapbuf_size3 mux_right_track_224 (
		.in({chany_top_in[111], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_311_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_311_sram_inv[0:1]),
		.out(chanx_right_out[112]));

	mux_tree_tapbuf_size3 mux_right_track_226 (
		.in({chany_top_in[112], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_312_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_312_sram_inv[0:1]),
		.out(chanx_right_out[113]));

	mux_tree_tapbuf_size3 mux_right_track_228 (
		.in({chany_top_in[113], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_313_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_313_sram_inv[0:1]),
		.out(chanx_right_out[114]));

	mux_tree_tapbuf_size3 mux_right_track_234 (
		.in({chany_top_in[116], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_314_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_314_sram_inv[0:1]),
		.out(chanx_right_out[117]));

	mux_tree_tapbuf_size3 mux_right_track_236 (
		.in({chany_top_in[117], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_315_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_315_sram_inv[0:1]),
		.out(chanx_right_out[118]));

	mux_tree_tapbuf_size3 mux_right_track_238 (
		.in({chany_top_in[118], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_316_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_316_sram_inv[0:1]),
		.out(chanx_right_out[119]));

	mux_tree_tapbuf_size3 mux_right_track_240 (
		.in({chany_top_in[119], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_317_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_317_sram_inv[0:1]),
		.out(chanx_right_out[120]));

	mux_tree_tapbuf_size3 mux_right_track_242 (
		.in({chany_top_in[120], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_318_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_318_sram_inv[0:1]),
		.out(chanx_right_out[121]));

	mux_tree_tapbuf_size3 mux_right_track_244 (
		.in({chany_top_in[121], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_319_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_319_sram_inv[0:1]),
		.out(chanx_right_out[122]));

	mux_tree_tapbuf_size3 mux_right_track_246 (
		.in({chany_top_in[122], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_320_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_320_sram_inv[0:1]),
		.out(chanx_right_out[123]));

	mux_tree_tapbuf_size3 mux_right_track_252 (
		.in({chany_top_in[125], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_321_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_321_sram_inv[0:1]),
		.out(chanx_right_out[126]));

	mux_tree_tapbuf_size3 mux_right_track_254 (
		.in({chany_top_in[126], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_322_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_322_sram_inv[0:1]),
		.out(chanx_right_out[127]));

	mux_tree_tapbuf_size3 mux_right_track_256 (
		.in({chany_top_in[127], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_323_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_323_sram_inv[0:1]),
		.out(chanx_right_out[128]));

	mux_tree_tapbuf_size3 mux_right_track_258 (
		.in({chany_top_in[128], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_324_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_324_sram_inv[0:1]),
		.out(chanx_right_out[129]));

	mux_tree_tapbuf_size3 mux_right_track_260 (
		.in({chany_top_in[129], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_325_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_325_sram_inv[0:1]),
		.out(chanx_right_out[130]));

	mux_tree_tapbuf_size3 mux_right_track_262 (
		.in({chany_top_in[130], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_326_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_326_sram_inv[0:1]),
		.out(chanx_right_out[131]));

	mux_tree_tapbuf_size3 mux_right_track_264 (
		.in({chany_top_in[131], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_327_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_327_sram_inv[0:1]),
		.out(chanx_right_out[132]));

	mux_tree_tapbuf_size3 mux_right_track_270 (
		.in({chany_top_in[134], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_328_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_328_sram_inv[0:1]),
		.out(chanx_right_out[135]));

	mux_tree_tapbuf_size3 mux_right_track_272 (
		.in({chany_top_in[135], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_329_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_329_sram_inv[0:1]),
		.out(chanx_right_out[136]));

	mux_tree_tapbuf_size3 mux_right_track_274 (
		.in({chany_top_in[136], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_330_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_330_sram_inv[0:1]),
		.out(chanx_right_out[137]));

	mux_tree_tapbuf_size3 mux_right_track_276 (
		.in({chany_top_in[137], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_331_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_331_sram_inv[0:1]),
		.out(chanx_right_out[138]));

	mux_tree_tapbuf_size3 mux_right_track_278 (
		.in({chany_top_in[138], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_332_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_332_sram_inv[0:1]),
		.out(chanx_right_out[139]));

	mux_tree_tapbuf_size3 mux_right_track_280 (
		.in({chany_top_in[139], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_333_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_333_sram_inv[0:1]),
		.out(chanx_right_out[140]));

	mux_tree_tapbuf_size3 mux_right_track_282 (
		.in({chany_top_in[140], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_334_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_334_sram_inv[0:1]),
		.out(chanx_right_out[141]));

	mux_tree_tapbuf_size3 mux_right_track_288 (
		.in({chany_top_in[143], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_335_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_335_sram_inv[0:1]),
		.out(chanx_right_out[144]));

	mux_tree_tapbuf_size3 mux_right_track_290 (
		.in({chany_top_in[144], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_336_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_336_sram_inv[0:1]),
		.out(chanx_right_out[145]));

	mux_tree_tapbuf_size3 mux_right_track_292 (
		.in({chany_top_in[145], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_337_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_337_sram_inv[0:1]),
		.out(chanx_right_out[146]));

	mux_tree_tapbuf_size3 mux_right_track_294 (
		.in({chany_top_in[146], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_338_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_338_sram_inv[0:1]),
		.out(chanx_right_out[147]));

	mux_tree_tapbuf_size3 mux_right_track_296 (
		.in({chany_top_in[147], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_339_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_339_sram_inv[0:1]),
		.out(chanx_right_out[148]));

	mux_tree_tapbuf_size3 mux_right_track_298 (
		.in({chany_top_in[148], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_340_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_340_sram_inv[0:1]),
		.out(chanx_right_out[149]));

	mux_tree_tapbuf_size3 mux_right_track_300 (
		.in({chany_top_in[149], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_341_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_341_sram_inv[0:1]),
		.out(chanx_right_out[150]));

	mux_tree_tapbuf_size3 mux_right_track_306 (
		.in({chany_top_in[152], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_342_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_342_sram_inv[0:1]),
		.out(chanx_right_out[153]));

	mux_tree_tapbuf_size3 mux_right_track_308 (
		.in({chany_top_in[153], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_343_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_343_sram_inv[0:1]),
		.out(chanx_right_out[154]));

	mux_tree_tapbuf_size3 mux_right_track_310 (
		.in({chany_top_in[154], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_344_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_344_sram_inv[0:1]),
		.out(chanx_right_out[155]));

	mux_tree_tapbuf_size3 mux_right_track_312 (
		.in({chany_top_in[155], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_345_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_345_sram_inv[0:1]),
		.out(chanx_right_out[156]));

	mux_tree_tapbuf_size3 mux_right_track_314 (
		.in({chany_top_in[156], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_346_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_346_sram_inv[0:1]),
		.out(chanx_right_out[157]));

	mux_tree_tapbuf_size3 mux_right_track_316 (
		.in({chany_top_in[157], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_347_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_347_sram_inv[0:1]),
		.out(chanx_right_out[158]));

	mux_tree_tapbuf_size3 mux_right_track_318 (
		.in({chany_top_in[158], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_348_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_348_sram_inv[0:1]),
		.out(chanx_right_out[159]));

	mux_tree_tapbuf_size3 mux_right_track_324 (
		.in({chany_top_in[161], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_349_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_349_sram_inv[0:1]),
		.out(chanx_right_out[162]));

	mux_tree_tapbuf_size3 mux_right_track_326 (
		.in({chany_top_in[162], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_350_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_350_sram_inv[0:1]),
		.out(chanx_right_out[163]));

	mux_tree_tapbuf_size3 mux_right_track_328 (
		.in({chany_top_in[163], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_351_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_351_sram_inv[0:1]),
		.out(chanx_right_out[164]));

	mux_tree_tapbuf_size3 mux_right_track_330 (
		.in({chany_top_in[164], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_352_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_352_sram_inv[0:1]),
		.out(chanx_right_out[165]));

	mux_tree_tapbuf_size3 mux_right_track_332 (
		.in({chany_top_in[165], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_353_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_353_sram_inv[0:1]),
		.out(chanx_right_out[166]));

	mux_tree_tapbuf_size3 mux_right_track_334 (
		.in({chany_top_in[166], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_354_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_354_sram_inv[0:1]),
		.out(chanx_right_out[167]));

	mux_tree_tapbuf_size3 mux_right_track_336 (
		.in({chany_top_in[167], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_355_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_355_sram_inv[0:1]),
		.out(chanx_right_out[168]));

	mux_tree_tapbuf_size3 mux_right_track_342 (
		.in({chany_top_in[170], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_356_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_356_sram_inv[0:1]),
		.out(chanx_right_out[171]));

	mux_tree_tapbuf_size3 mux_right_track_344 (
		.in({chany_top_in[171], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_357_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_357_sram_inv[0:1]),
		.out(chanx_right_out[172]));

	mux_tree_tapbuf_size3 mux_right_track_346 (
		.in({chany_top_in[172], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_358_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_358_sram_inv[0:1]),
		.out(chanx_right_out[173]));

	mux_tree_tapbuf_size3 mux_right_track_348 (
		.in({chany_top_in[173], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_359_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_359_sram_inv[0:1]),
		.out(chanx_right_out[174]));

	mux_tree_tapbuf_size3 mux_right_track_350 (
		.in({chany_top_in[174], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_360_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_360_sram_inv[0:1]),
		.out(chanx_right_out[175]));

	mux_tree_tapbuf_size3 mux_right_track_352 (
		.in({chany_top_in[175], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_361_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_361_sram_inv[0:1]),
		.out(chanx_right_out[176]));

	mux_tree_tapbuf_size3 mux_right_track_354 (
		.in({chany_top_in[176], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_362_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_362_sram_inv[0:1]),
		.out(chanx_right_out[177]));

	mux_tree_tapbuf_size3 mux_right_track_360 (
		.in({chany_top_in[179], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_363_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_363_sram_inv[0:1]),
		.out(chanx_right_out[180]));

	mux_tree_tapbuf_size3 mux_right_track_362 (
		.in({chany_top_in[180], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_364_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_364_sram_inv[0:1]),
		.out(chanx_right_out[181]));

	mux_tree_tapbuf_size3 mux_right_track_364 (
		.in({chany_top_in[181], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_365_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_365_sram_inv[0:1]),
		.out(chanx_right_out[182]));

	mux_tree_tapbuf_size3 mux_right_track_366 (
		.in({chany_top_in[182], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_366_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_366_sram_inv[0:1]),
		.out(chanx_right_out[183]));

	mux_tree_tapbuf_size3 mux_right_track_368 (
		.in({chany_top_in[183], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_367_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_367_sram_inv[0:1]),
		.out(chanx_right_out[184]));

	mux_tree_tapbuf_size3 mux_right_track_370 (
		.in({chany_top_in[184], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_368_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_368_sram_inv[0:1]),
		.out(chanx_right_out[185]));

	mux_tree_tapbuf_size3 mux_right_track_372 (
		.in({chany_top_in[185], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_369_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_369_sram_inv[0:1]),
		.out(chanx_right_out[186]));

	mux_tree_tapbuf_size3 mux_right_track_378 (
		.in({chany_top_in[188], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_370_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_370_sram_inv[0:1]),
		.out(chanx_right_out[189]));

	mux_tree_tapbuf_size3 mux_right_track_380 (
		.in({chany_top_in[189], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_371_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_371_sram_inv[0:1]),
		.out(chanx_right_out[190]));

	mux_tree_tapbuf_size3 mux_right_track_382 (
		.in({chany_top_in[190], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_372_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_372_sram_inv[0:1]),
		.out(chanx_right_out[191]));

	mux_tree_tapbuf_size3 mux_right_track_384 (
		.in({chany_top_in[191], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_373_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_373_sram_inv[0:1]),
		.out(chanx_right_out[192]));

	mux_tree_tapbuf_size3 mux_right_track_386 (
		.in({chany_top_in[192], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_374_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_374_sram_inv[0:1]),
		.out(chanx_right_out[193]));

	mux_tree_tapbuf_size3 mux_right_track_388 (
		.in({chany_top_in[193], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_375_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_375_sram_inv[0:1]),
		.out(chanx_right_out[194]));

	mux_tree_tapbuf_size3 mux_right_track_390 (
		.in({chany_top_in[194], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_376_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_376_sram_inv[0:1]),
		.out(chanx_right_out[195]));

	mux_tree_tapbuf_size3 mux_right_track_396 (
		.in({chany_top_in[197], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_377_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_377_sram_inv[0:1]),
		.out(chanx_right_out[198]));

	mux_tree_tapbuf_size3 mux_right_track_398 (
		.in({chany_top_in[198], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_378_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_378_sram_inv[0:1]),
		.out(chanx_right_out[199]));

	mux_tree_tapbuf_size3 mux_right_track_400 (
		.in({chany_top_in[199], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_379_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_379_sram_inv[0:1]),
		.out(chanx_right_out[200]));

	mux_tree_tapbuf_size3 mux_right_track_402 (
		.in({chany_top_in[200], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_380_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_380_sram_inv[0:1]),
		.out(chanx_right_out[201]));

	mux_tree_tapbuf_size3 mux_right_track_404 (
		.in({chany_top_in[201], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_381_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_381_sram_inv[0:1]),
		.out(chanx_right_out[202]));

	mux_tree_tapbuf_size3 mux_right_track_406 (
		.in({chany_top_in[202], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_382_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_382_sram_inv[0:1]),
		.out(chanx_right_out[203]));

	mux_tree_tapbuf_size3 mux_right_track_408 (
		.in({chany_top_in[203], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_383_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_383_sram_inv[0:1]),
		.out(chanx_right_out[204]));

	mux_tree_tapbuf_size3 mux_right_track_414 (
		.in({chany_top_in[206], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_384_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_384_sram_inv[0:1]),
		.out(chanx_right_out[207]));

	mux_tree_tapbuf_size3 mux_right_track_416 (
		.in({chany_top_in[207], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_385_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_385_sram_inv[0:1]),
		.out(chanx_right_out[208]));

	mux_tree_tapbuf_size3 mux_right_track_418 (
		.in({chany_top_in[208], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_386_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_386_sram_inv[0:1]),
		.out(chanx_right_out[209]));

	mux_tree_tapbuf_size3 mux_right_track_420 (
		.in({chany_top_in[209], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_387_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_387_sram_inv[0:1]),
		.out(chanx_right_out[210]));

	mux_tree_tapbuf_size3 mux_right_track_422 (
		.in({chany_top_in[210], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_388_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_388_sram_inv[0:1]),
		.out(chanx_right_out[211]));

	mux_tree_tapbuf_size3 mux_right_track_424 (
		.in({chany_top_in[211], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_389_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_389_sram_inv[0:1]),
		.out(chanx_right_out[212]));

	mux_tree_tapbuf_size3 mux_right_track_426 (
		.in({chany_top_in[212], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_390_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_390_sram_inv[0:1]),
		.out(chanx_right_out[213]));

	mux_tree_tapbuf_size3 mux_right_track_432 (
		.in({chany_top_in[215], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_391_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_391_sram_inv[0:1]),
		.out(chanx_right_out[216]));

	mux_tree_tapbuf_size3 mux_right_track_434 (
		.in({chany_top_in[216], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_392_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_392_sram_inv[0:1]),
		.out(chanx_right_out[217]));

	mux_tree_tapbuf_size3 mux_right_track_436 (
		.in({chany_top_in[217], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_393_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_393_sram_inv[0:1]),
		.out(chanx_right_out[218]));

	mux_tree_tapbuf_size3 mux_right_track_438 (
		.in({chany_top_in[218], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_394_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_394_sram_inv[0:1]),
		.out(chanx_right_out[219]));

	mux_tree_tapbuf_size3 mux_right_track_440 (
		.in({chany_top_in[219], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_395_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_395_sram_inv[0:1]),
		.out(chanx_right_out[220]));

	mux_tree_tapbuf_size3 mux_right_track_442 (
		.in({chany_top_in[220], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_396_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_396_sram_inv[0:1]),
		.out(chanx_right_out[221]));

	mux_tree_tapbuf_size3 mux_right_track_444 (
		.in({chany_top_in[221], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_397_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_397_sram_inv[0:1]),
		.out(chanx_right_out[222]));

	mux_tree_tapbuf_size3 mux_right_track_450 (
		.in({chany_top_in[224], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_398_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_398_sram_inv[0:1]),
		.out(chanx_right_out[225]));

	mux_tree_tapbuf_size3 mux_right_track_452 (
		.in({chany_top_in[225], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_399_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_399_sram_inv[0:1]),
		.out(chanx_right_out[226]));

	mux_tree_tapbuf_size3 mux_right_track_454 (
		.in({chany_top_in[226], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_400_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_400_sram_inv[0:1]),
		.out(chanx_right_out[227]));

	mux_tree_tapbuf_size3 mux_right_track_456 (
		.in({chany_top_in[227], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_401_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_401_sram_inv[0:1]),
		.out(chanx_right_out[228]));

	mux_tree_tapbuf_size3 mux_right_track_458 (
		.in({chany_top_in[228], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_402_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_402_sram_inv[0:1]),
		.out(chanx_right_out[229]));

	mux_tree_tapbuf_size3 mux_right_track_460 (
		.in({chany_top_in[229], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_403_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_403_sram_inv[0:1]),
		.out(chanx_right_out[230]));

	mux_tree_tapbuf_size3 mux_right_track_462 (
		.in({chany_top_in[230], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_404_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_404_sram_inv[0:1]),
		.out(chanx_right_out[231]));

	mux_tree_tapbuf_size3 mux_right_track_468 (
		.in({chany_top_in[233], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_405_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_405_sram_inv[0:1]),
		.out(chanx_right_out[234]));

	mux_tree_tapbuf_size3 mux_right_track_470 (
		.in({chany_top_in[234], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_406_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_406_sram_inv[0:1]),
		.out(chanx_right_out[235]));

	mux_tree_tapbuf_size3 mux_right_track_472 (
		.in({chany_top_in[235], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_407_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_407_sram_inv[0:1]),
		.out(chanx_right_out[236]));

	mux_tree_tapbuf_size3 mux_right_track_474 (
		.in({chany_top_in[236], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_408_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_408_sram_inv[0:1]),
		.out(chanx_right_out[237]));

	mux_tree_tapbuf_size3 mux_right_track_476 (
		.in({chany_top_in[237], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_409_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_409_sram_inv[0:1]),
		.out(chanx_right_out[238]));

	mux_tree_tapbuf_size3 mux_right_track_478 (
		.in({chany_top_in[238], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_410_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_410_sram_inv[0:1]),
		.out(chanx_right_out[239]));

	mux_tree_tapbuf_size3 mux_right_track_480 (
		.in({chany_top_in[239], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_411_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_411_sram_inv[0:1]),
		.out(chanx_right_out[240]));

	mux_tree_tapbuf_size3 mux_right_track_486 (
		.in({chany_top_in[242], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_412_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_412_sram_inv[0:1]),
		.out(chanx_right_out[243]));

	mux_tree_tapbuf_size3 mux_right_track_488 (
		.in({chany_top_in[243], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_413_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_413_sram_inv[0:1]),
		.out(chanx_right_out[244]));

	mux_tree_tapbuf_size3 mux_right_track_490 (
		.in({chany_top_in[244], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_414_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_414_sram_inv[0:1]),
		.out(chanx_right_out[245]));

	mux_tree_tapbuf_size3 mux_right_track_492 (
		.in({chany_top_in[245], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_415_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_415_sram_inv[0:1]),
		.out(chanx_right_out[246]));

	mux_tree_tapbuf_size3 mux_right_track_494 (
		.in({chany_top_in[246], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_416_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_416_sram_inv[0:1]),
		.out(chanx_right_out[247]));

	mux_tree_tapbuf_size3 mux_right_track_496 (
		.in({chany_top_in[247], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_417_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_417_sram_inv[0:1]),
		.out(chanx_right_out[248]));

	mux_tree_tapbuf_size3 mux_right_track_498 (
		.in({chany_top_in[248], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_418_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_418_sram_inv[0:1]),
		.out(chanx_right_out[249]));

	mux_tree_tapbuf_size3 mux_right_track_504 (
		.in({chany_top_in[251], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_419_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_419_sram_inv[0:1]),
		.out(chanx_right_out[252]));

	mux_tree_tapbuf_size3 mux_right_track_506 (
		.in({chany_top_in[252], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_420_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_420_sram_inv[0:1]),
		.out(chanx_right_out[253]));

	mux_tree_tapbuf_size3 mux_right_track_508 (
		.in({chany_top_in[253], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_421_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_421_sram_inv[0:1]),
		.out(chanx_right_out[254]));

	mux_tree_tapbuf_size3 mux_right_track_510 (
		.in({chany_top_in[254], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_422_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_422_sram_inv[0:1]),
		.out(chanx_right_out[255]));

	mux_tree_tapbuf_size3 mux_right_track_512 (
		.in({chany_top_in[255], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_423_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_423_sram_inv[0:1]),
		.out(chanx_right_out[256]));

	mux_tree_tapbuf_size3 mux_right_track_514 (
		.in({chany_top_in[256], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_424_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_424_sram_inv[0:1]),
		.out(chanx_right_out[257]));

	mux_tree_tapbuf_size3 mux_right_track_516 (
		.in({chany_top_in[257], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_425_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_425_sram_inv[0:1]),
		.out(chanx_right_out[258]));

	mux_tree_tapbuf_size3 mux_right_track_522 (
		.in({chany_top_in[260], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_426_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_426_sram_inv[0:1]),
		.out(chanx_right_out[261]));

	mux_tree_tapbuf_size3 mux_right_track_524 (
		.in({chany_top_in[261], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_427_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_427_sram_inv[0:1]),
		.out(chanx_right_out[262]));

	mux_tree_tapbuf_size3 mux_right_track_526 (
		.in({chany_top_in[262], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_428_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_428_sram_inv[0:1]),
		.out(chanx_right_out[263]));

	mux_tree_tapbuf_size3 mux_right_track_528 (
		.in({chany_top_in[263], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_429_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_429_sram_inv[0:1]),
		.out(chanx_right_out[264]));

	mux_tree_tapbuf_size3 mux_right_track_530 (
		.in({chany_top_in[264], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_430_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_430_sram_inv[0:1]),
		.out(chanx_right_out[265]));

	mux_tree_tapbuf_size3 mux_right_track_532 (
		.in({chany_top_in[265], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_431_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_431_sram_inv[0:1]),
		.out(chanx_right_out[266]));

	mux_tree_tapbuf_size3 mux_right_track_534 (
		.in({chany_top_in[266], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_432_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_432_sram_inv[0:1]),
		.out(chanx_right_out[267]));

	mux_tree_tapbuf_size3 mux_right_track_540 (
		.in({chany_top_in[269], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_433_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_433_sram_inv[0:1]),
		.out(chanx_right_out[270]));

	mux_tree_tapbuf_size3 mux_right_track_542 (
		.in({chany_top_in[270], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_434_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_434_sram_inv[0:1]),
		.out(chanx_right_out[271]));

	mux_tree_tapbuf_size3 mux_right_track_544 (
		.in({chany_top_in[271], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_435_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_435_sram_inv[0:1]),
		.out(chanx_right_out[272]));

	mux_tree_tapbuf_size3 mux_right_track_546 (
		.in({chany_top_in[272], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_436_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_436_sram_inv[0:1]),
		.out(chanx_right_out[273]));

	mux_tree_tapbuf_size3 mux_right_track_548 (
		.in({chany_top_in[273], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_437_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_437_sram_inv[0:1]),
		.out(chanx_right_out[274]));

	mux_tree_tapbuf_size3 mux_right_track_550 (
		.in({chany_top_in[274], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_438_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_438_sram_inv[0:1]),
		.out(chanx_right_out[275]));

	mux_tree_tapbuf_size3 mux_right_track_552 (
		.in({chany_top_in[275], right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_439_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_439_sram_inv[0:1]),
		.out(chanx_right_out[276]));

	mux_tree_tapbuf_size3 mux_right_track_558 (
		.in({chany_top_in[278], right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_440_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_440_sram_inv[0:1]),
		.out(chanx_right_out[279]));

	mux_tree_tapbuf_size3 mux_right_track_560 (
		.in({chany_top_in[279], right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_441_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_441_sram_inv[0:1]),
		.out(chanx_right_out[280]));

	mux_tree_tapbuf_size3 mux_right_track_562 (
		.in({chany_top_in[280], right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_442_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_442_sram_inv[0:1]),
		.out(chanx_right_out[281]));

	mux_tree_tapbuf_size3 mux_right_track_564 (
		.in({chany_top_in[281], right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_443_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_443_sram_inv[0:1]),
		.out(chanx_right_out[282]));

	mux_tree_tapbuf_size3 mux_right_track_566 (
		.in({chany_top_in[282], right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_444_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_444_sram_inv[0:1]),
		.out(chanx_right_out[283]));

	mux_tree_tapbuf_size3 mux_right_track_568 (
		.in({chany_top_in[283], right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_, right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size3_445_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size3_445_sram_inv[0:1]),
		.out(chanx_right_out[284]));

	mux_tree_tapbuf_size3_mem mem_top_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_0_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_1_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_2_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_3_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_4_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_5_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_6_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_7_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_8_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_9_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_10_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_11_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_12_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_13_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_14_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_15_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_16_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_17_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_18_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_19_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_20_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_21_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_22_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_23_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_24_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_25_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_26_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_27_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_28_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_29_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_30_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_31_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_32_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_33_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_34_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_35_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_36_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_37_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_38_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_39_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_40_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_41_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_42_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_43_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_44_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_45_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_46_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_47_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_48_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_49_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_50_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_51_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_52_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_53_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_54_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_55_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_56_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_57_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_58_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_59_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_60_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_61_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_62_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_63_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_64_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_65_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_66_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_67_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_68_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_69_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_70_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_71_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_72_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_73_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_74_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_75_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_76_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_77_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_78_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_79_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_80_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_81_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_82_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_83_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_84_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_85_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_86_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_87_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_88_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_89_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_90_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_91_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_92_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_93_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_94_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_95_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_96_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_97_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_98_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_99_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_100_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_101_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_102_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_103_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_104_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_105_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_106_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_107_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_108_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_109_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_110_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_111_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_112_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_113_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_114_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_115_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_116_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_117_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_118_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_119_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_120_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_120_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_120_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_121_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_121_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_121_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_122_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_122_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_122_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_123_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_123_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_123_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_124_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_124_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_124_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_125_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_125_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_126_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_126_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_126_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_127_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_127_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_127_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_128_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_128_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_128_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_129_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_129_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_129_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_130_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_130_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_130_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_131_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_131_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_131_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_132_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_132_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_133_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_133_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_133_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_134_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_134_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_134_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_135_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_135_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_135_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_136_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_136_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_136_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_137_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_137_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_137_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_138_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_138_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_138_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_139_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_139_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_140_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_140_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_140_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_141_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_141_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_141_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_142_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_142_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_142_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_143_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_143_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_143_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_144_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_144_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_144_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_145_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_145_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_145_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_146_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_146_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_378 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_147_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_147_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_380 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_147_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_148_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_148_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_382 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_148_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_149_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_149_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_149_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_150_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_150_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_386 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_150_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_151_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_151_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_388 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_151_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_152_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_152_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_390 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_152_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_153_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_153_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_396 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_154_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_154_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_398 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_154_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_155_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_155_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_155_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_156_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_156_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_402 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_156_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_157_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_157_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_404 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_157_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_158_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_158_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_406 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_158_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_159_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_159_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_159_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_160_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_160_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_414 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_161_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_161_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_161_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_162_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_162_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_418 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_162_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_163_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_163_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_420 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_163_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_164_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_164_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_422 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_164_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_165_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_165_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_165_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_166_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_166_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_426 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_166_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_167_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_167_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_168_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_168_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_434 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_168_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_169_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_169_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_436 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_169_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_170_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_170_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_438 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_170_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_171_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_171_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_171_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_171_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_172_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_172_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_172_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_442 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_172_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_173_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_173_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_173_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_444 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_173_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_174_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_174_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_174_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_450 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_175_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_175_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_175_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_452 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_175_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_176_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_176_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_176_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_454 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_176_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_177_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_177_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_177_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_177_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_178_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_178_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_178_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_458 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_178_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_179_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_179_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_179_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_460 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_179_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_180_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_180_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_180_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_462 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_180_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_181_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_181_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_181_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_468 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_182_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_182_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_182_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_470 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_182_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_183_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_183_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_183_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_183_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_184_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_184_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_184_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_474 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_184_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_185_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_185_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_185_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_476 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_185_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_186_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_186_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_186_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_478 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_186_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_187_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_187_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_187_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_187_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_188_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_188_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_188_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_486 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_189_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_189_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_189_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_189_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_190_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_190_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_190_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_490 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_190_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_191_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_191_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_191_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_492 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_191_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_192_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_192_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_192_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_494 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_192_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_193_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_193_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_193_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_193_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_194_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_194_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_194_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_498 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_194_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_195_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_195_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_195_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_196_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_196_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_196_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_506 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_196_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_197_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_197_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_197_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_508 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_197_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_198_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_198_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_198_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_510 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_198_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_199_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_199_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_199_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_199_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_200_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_200_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_200_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_514 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_200_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_201_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_201_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_201_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_516 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_201_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_202_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_202_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_202_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_522 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_203_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_203_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_203_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_524 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_203_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_204_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_204_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_204_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_526 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_204_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_205_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_205_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_205_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_205_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_206_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_206_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_206_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_530 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_206_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_207_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_207_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_207_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_532 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_207_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_208_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_208_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_208_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_534 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_208_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_209_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_209_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_209_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_540 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_210_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_210_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_210_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_542 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_210_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_211_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_211_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_211_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_211_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_212_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_212_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_212_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_546 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_212_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_213_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_213_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_213_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_548 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_213_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_214_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_214_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_214_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_550 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_214_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_215_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_215_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_215_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_215_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_216_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_216_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_216_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_558 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_217_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_217_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_217_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_217_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_218_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_218_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_218_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_562 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_218_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_219_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_219_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_219_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_564 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_219_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_220_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_220_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_220_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_566 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_220_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_221_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_221_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_221_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_top_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_221_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_222_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_222_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_222_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_223_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_223_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_223_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_223_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_224_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_224_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_224_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_224_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_225_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_225_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_225_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_225_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_226_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_226_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_226_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_226_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_227_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_227_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_227_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_227_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_228_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_228_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_228_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_228_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_229_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_229_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_229_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_229_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_230_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_230_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_230_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size4_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_231_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_231_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_231_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_231_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_232_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_232_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_232_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_232_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_233_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_233_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_233_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_233_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_234_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_234_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_234_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_234_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_235_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_235_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_235_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_235_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_236_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_236_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_236_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_237_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_237_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_237_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_237_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_238_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_238_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_238_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_238_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_239_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_239_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_239_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_239_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_240_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_240_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_240_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_240_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_241_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_241_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_241_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_241_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_242_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_242_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_242_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_242_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_243_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_243_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_243_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_244_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_244_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_244_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_244_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_245_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_245_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_245_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_245_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_246_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_246_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_246_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_246_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_247_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_247_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_247_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_247_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_248_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_248_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_248_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_248_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_249_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_249_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_249_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_249_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_250_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_250_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_250_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_251_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_251_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_251_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_251_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_252_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_252_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_252_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_252_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_253_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_253_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_253_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_253_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_254_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_254_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_254_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_254_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_255_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_255_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_255_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_255_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_256_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_256_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_256_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_256_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_257_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_257_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_257_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_258_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_258_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_258_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_258_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_259_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_259_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_259_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_259_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_260_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_260_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_260_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_260_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_261_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_261_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_261_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_261_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_262_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_262_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_262_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_262_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_263_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_263_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_263_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_263_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_264_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_264_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_264_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_265_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_265_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_265_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_265_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_266_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_266_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_266_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_266_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_267_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_267_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_267_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_267_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_268_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_268_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_268_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_268_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_269_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_269_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_269_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_269_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_270_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_270_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_270_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_270_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_271_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_271_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_271_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_272_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_272_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_272_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_272_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_273_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_273_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_273_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_273_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_274_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_274_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_274_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_274_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_275_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_275_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_275_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_275_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_276_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_276_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_276_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_276_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_277_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_277_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_277_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_277_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_278_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_278_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_278_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_279_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_279_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_279_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_146 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_279_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_280_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_280_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_280_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_148 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_280_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_281_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_281_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_281_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_150 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_281_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_282_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_282_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_282_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_152 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_282_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_283_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_283_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_283_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_154 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_283_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_284_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_284_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_284_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_156 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_284_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_285_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_285_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_285_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_162 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_286_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_286_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_286_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_164 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_286_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_287_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_287_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_287_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_166 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_287_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_288_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_288_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_288_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_168 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_288_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_289_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_289_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_289_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_170 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_289_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_290_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_290_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_290_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_172 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_290_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_291_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_291_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_291_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_174 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_291_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_292_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_292_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_292_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_180 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_293_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_293_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_293_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_182 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_293_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_294_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_294_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_294_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_184 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_294_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_295_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_295_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_295_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_186 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_295_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_296_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_296_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_296_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_188 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_296_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_297_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_297_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_297_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_190 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_297_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_298_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_298_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_298_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_192 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_298_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_299_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_299_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_299_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_198 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_300_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_300_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_300_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_200 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_300_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_301_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_301_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_301_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_202 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_301_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_302_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_302_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_302_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_204 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_302_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_303_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_303_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_303_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_206 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_303_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_304_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_304_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_304_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_208 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_304_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_305_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_305_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_305_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_210 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_305_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_306_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_306_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_306_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_216 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_307_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_307_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_307_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_218 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_307_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_308_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_308_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_308_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_220 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_308_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_309_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_309_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_309_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_222 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_309_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_310_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_310_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_310_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_224 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_310_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_311_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_311_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_311_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_226 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_311_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_312_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_312_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_312_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_228 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_312_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_313_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_313_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_313_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_234 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_314_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_314_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_314_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_236 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_314_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_315_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_315_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_315_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_238 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_315_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_316_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_316_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_316_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_240 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_316_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_317_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_317_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_317_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_242 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_317_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_318_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_318_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_318_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_244 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_318_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_319_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_319_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_319_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_246 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_319_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_320_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_320_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_320_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_252 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_321_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_321_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_321_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_254 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_321_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_322_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_322_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_322_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_256 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_322_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_323_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_323_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_323_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_258 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_323_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_324_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_324_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_324_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_260 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_324_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_325_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_325_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_325_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_262 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_325_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_326_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_326_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_326_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_264 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_326_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_327_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_327_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_327_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_270 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_328_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_328_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_328_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_272 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_328_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_329_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_329_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_329_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_274 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_329_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_330_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_330_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_330_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_276 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_330_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_331_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_331_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_331_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_278 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_331_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_332_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_332_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_332_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_280 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_332_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_333_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_333_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_333_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_282 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_333_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_334_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_334_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_334_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_288 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_335_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_335_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_335_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_290 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_335_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_336_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_336_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_336_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_292 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_336_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_337_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_337_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_337_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_294 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_337_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_338_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_338_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_338_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_296 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_338_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_339_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_339_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_339_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_298 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_339_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_340_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_340_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_340_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_300 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_340_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_341_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_341_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_341_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_306 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_342_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_342_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_342_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_308 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_342_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_343_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_343_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_343_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_310 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_343_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_344_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_344_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_344_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_312 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_344_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_345_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_345_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_345_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_314 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_345_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_346_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_346_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_346_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_316 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_346_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_347_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_347_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_347_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_318 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_347_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_348_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_348_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_348_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_324 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_349_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_349_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_349_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_326 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_349_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_350_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_350_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_350_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_328 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_350_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_351_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_351_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_351_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_330 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_351_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_352_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_352_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_352_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_332 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_352_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_353_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_353_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_353_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_334 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_353_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_354_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_354_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_354_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_336 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_354_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_355_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_355_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_355_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_342 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_356_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_356_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_356_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_344 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_356_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_357_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_357_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_357_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_346 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_357_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_358_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_358_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_358_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_348 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_358_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_359_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_359_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_359_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_350 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_359_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_360_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_360_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_360_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_352 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_360_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_361_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_361_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_361_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_354 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_361_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_362_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_362_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_362_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_360 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_363_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_363_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_363_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_362 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_363_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_364_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_364_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_364_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_364 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_364_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_365_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_365_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_365_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_366 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_365_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_366_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_366_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_366_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_368 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_366_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_367_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_367_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_367_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_370 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_367_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_368_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_368_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_368_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_372 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_368_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_369_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_369_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_369_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_378 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_370_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_370_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_370_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_380 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_370_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_371_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_371_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_371_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_382 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_371_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_372_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_372_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_372_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_384 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_372_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_373_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_373_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_373_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_386 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_373_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_374_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_374_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_374_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_388 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_374_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_375_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_375_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_375_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_390 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_375_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_376_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_376_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_376_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_396 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_377_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_377_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_377_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_398 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_377_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_378_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_378_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_378_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_400 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_378_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_379_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_379_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_379_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_402 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_379_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_380_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_380_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_380_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_404 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_380_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_381_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_381_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_381_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_406 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_381_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_382_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_382_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_382_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_408 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_382_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_383_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_383_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_383_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_414 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_384_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_384_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_384_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_416 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_384_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_385_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_385_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_385_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_418 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_385_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_386_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_386_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_386_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_420 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_386_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_387_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_387_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_387_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_422 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_387_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_388_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_388_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_388_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_424 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_388_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_389_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_389_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_389_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_426 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_389_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_390_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_390_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_390_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_432 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_391_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_391_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_391_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_434 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_391_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_392_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_392_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_392_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_436 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_392_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_393_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_393_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_393_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_438 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_393_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_394_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_394_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_394_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_440 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_394_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_395_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_395_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_395_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_442 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_395_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_396_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_396_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_396_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_444 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_396_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_397_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_397_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_397_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_450 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_398_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_398_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_398_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_452 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_398_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_399_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_399_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_399_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_454 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_399_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_400_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_400_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_400_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_456 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_400_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_401_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_401_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_401_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_458 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_401_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_402_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_402_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_402_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_460 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_402_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_403_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_403_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_403_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_462 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_403_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_404_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_404_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_404_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_468 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_405_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_405_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_405_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_470 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_405_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_406_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_406_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_406_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_472 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_406_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_407_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_407_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_407_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_474 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_407_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_408_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_408_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_408_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_476 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_408_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_409_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_409_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_409_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_478 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_409_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_410_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_410_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_410_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_480 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_410_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_411_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_411_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_411_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_486 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_412_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_412_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_412_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_488 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_412_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_413_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_413_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_413_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_490 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_413_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_414_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_414_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_414_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_492 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_414_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_415_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_415_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_415_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_494 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_415_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_416_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_416_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_416_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_496 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_416_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_417_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_417_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_417_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_498 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_417_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_418_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_418_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_418_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_504 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_419_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_419_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_419_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_506 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_419_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_420_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_420_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_420_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_508 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_420_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_421_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_421_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_421_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_510 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_421_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_422_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_422_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_422_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_512 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_422_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_423_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_423_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_423_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_514 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_423_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_424_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_424_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_424_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_516 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_424_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_425_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_425_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_425_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_522 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_426_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_426_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_426_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_524 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_426_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_427_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_427_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_427_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_526 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_427_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_428_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_428_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_428_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_528 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_428_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_429_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_429_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_429_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_530 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_429_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_430_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_430_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_430_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_532 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_430_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_431_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_431_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_431_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_534 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_431_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_432_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_432_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_432_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_540 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_433_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_433_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_433_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_542 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_433_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_434_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_434_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_434_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_544 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_434_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_435_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_435_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_435_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_546 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_435_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_436_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_436_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_436_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_548 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_436_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_437_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_437_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_437_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_550 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_437_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_438_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_438_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_438_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_552 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_438_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_439_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_439_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_439_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_558 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_440_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_440_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_440_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_560 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_440_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_441_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_441_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_441_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_562 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_441_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_442_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_442_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_442_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_564 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_442_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_443_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_443_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_443_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_566 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_443_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size3_mem_444_ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_444_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_444_sram_inv[0:1]));

	mux_tree_tapbuf_size3_mem mem_right_track_568 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_444_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size3_445_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size3_445_sram_inv[0:1]));

	mux_tree_tapbuf_size2 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[17]}),
		.sram(mux_tree_tapbuf_size2_0_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_0_sram_inv[0:1]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size2 mux_top_track_34 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[18]}),
		.sram(mux_tree_tapbuf_size2_1_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_1_sram_inv[0:1]),
		.out(chany_top_out[17]));

	mux_tree_tapbuf_size2 mux_top_track_50 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[26]}),
		.sram(mux_tree_tapbuf_size2_2_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_2_sram_inv[0:1]),
		.out(chany_top_out[25]));

	mux_tree_tapbuf_size2 mux_top_track_52 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[27]}),
		.sram(mux_tree_tapbuf_size2_3_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_3_sram_inv[0:1]),
		.out(chany_top_out[26]));

	mux_tree_tapbuf_size2 mux_top_track_68 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[35]}),
		.sram(mux_tree_tapbuf_size2_4_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_4_sram_inv[0:1]),
		.out(chany_top_out[34]));

	mux_tree_tapbuf_size2 mux_top_track_70 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[36]}),
		.sram(mux_tree_tapbuf_size2_5_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_5_sram_inv[0:1]),
		.out(chany_top_out[35]));

	mux_tree_tapbuf_size2 mux_top_track_86 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[44]}),
		.sram(mux_tree_tapbuf_size2_6_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_6_sram_inv[0:1]),
		.out(chany_top_out[43]));

	mux_tree_tapbuf_size2 mux_top_track_88 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[45]}),
		.sram(mux_tree_tapbuf_size2_7_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_7_sram_inv[0:1]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size2 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[53]}),
		.sram(mux_tree_tapbuf_size2_8_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_8_sram_inv[0:1]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size2 mux_top_track_106 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[54]}),
		.sram(mux_tree_tapbuf_size2_9_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_9_sram_inv[0:1]),
		.out(chany_top_out[53]));

	mux_tree_tapbuf_size2 mux_top_track_122 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[62]}),
		.sram(mux_tree_tapbuf_size2_10_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_10_sram_inv[0:1]),
		.out(chany_top_out[61]));

	mux_tree_tapbuf_size2 mux_top_track_124 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_size2_11_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_11_sram_inv[0:1]),
		.out(chany_top_out[62]));

	mux_tree_tapbuf_size2 mux_top_track_140 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_size2_12_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_12_sram_inv[0:1]),
		.out(chany_top_out[70]));

	mux_tree_tapbuf_size2 mux_top_track_142 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size2_13_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_13_sram_inv[0:1]),
		.out(chany_top_out[71]));

	mux_tree_tapbuf_size2 mux_top_track_158 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[80]}),
		.sram(mux_tree_tapbuf_size2_14_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_14_sram_inv[0:1]),
		.out(chany_top_out[79]));

	mux_tree_tapbuf_size2 mux_top_track_160 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[81]}),
		.sram(mux_tree_tapbuf_size2_15_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_15_sram_inv[0:1]),
		.out(chany_top_out[80]));

	mux_tree_tapbuf_size2 mux_top_track_176 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[89]}),
		.sram(mux_tree_tapbuf_size2_16_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_16_sram_inv[0:1]),
		.out(chany_top_out[88]));

	mux_tree_tapbuf_size2 mux_top_track_178 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[90]}),
		.sram(mux_tree_tapbuf_size2_17_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_17_sram_inv[0:1]),
		.out(chany_top_out[89]));

	mux_tree_tapbuf_size2 mux_top_track_194 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[98]}),
		.sram(mux_tree_tapbuf_size2_18_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_18_sram_inv[0:1]),
		.out(chany_top_out[97]));

	mux_tree_tapbuf_size2 mux_top_track_196 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[99]}),
		.sram(mux_tree_tapbuf_size2_19_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_19_sram_inv[0:1]),
		.out(chany_top_out[98]));

	mux_tree_tapbuf_size2 mux_top_track_212 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[107]}),
		.sram(mux_tree_tapbuf_size2_20_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_20_sram_inv[0:1]),
		.out(chany_top_out[106]));

	mux_tree_tapbuf_size2 mux_top_track_214 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[108]}),
		.sram(mux_tree_tapbuf_size2_21_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_21_sram_inv[0:1]),
		.out(chany_top_out[107]));

	mux_tree_tapbuf_size2 mux_top_track_230 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[116]}),
		.sram(mux_tree_tapbuf_size2_22_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_22_sram_inv[0:1]),
		.out(chany_top_out[115]));

	mux_tree_tapbuf_size2 mux_top_track_232 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[117]}),
		.sram(mux_tree_tapbuf_size2_23_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_23_sram_inv[0:1]),
		.out(chany_top_out[116]));

	mux_tree_tapbuf_size2 mux_top_track_248 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[125]}),
		.sram(mux_tree_tapbuf_size2_24_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_24_sram_inv[0:1]),
		.out(chany_top_out[124]));

	mux_tree_tapbuf_size2 mux_top_track_250 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[126]}),
		.sram(mux_tree_tapbuf_size2_25_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_25_sram_inv[0:1]),
		.out(chany_top_out[125]));

	mux_tree_tapbuf_size2 mux_top_track_266 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[134]}),
		.sram(mux_tree_tapbuf_size2_26_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_26_sram_inv[0:1]),
		.out(chany_top_out[133]));

	mux_tree_tapbuf_size2 mux_top_track_268 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[135]}),
		.sram(mux_tree_tapbuf_size2_27_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_27_sram_inv[0:1]),
		.out(chany_top_out[134]));

	mux_tree_tapbuf_size2 mux_top_track_284 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[143]}),
		.sram(mux_tree_tapbuf_size2_28_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_28_sram_inv[0:1]),
		.out(chany_top_out[142]));

	mux_tree_tapbuf_size2 mux_top_track_286 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[144]}),
		.sram(mux_tree_tapbuf_size2_29_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_29_sram_inv[0:1]),
		.out(chany_top_out[143]));

	mux_tree_tapbuf_size2 mux_top_track_302 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[152]}),
		.sram(mux_tree_tapbuf_size2_30_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_30_sram_inv[0:1]),
		.out(chany_top_out[151]));

	mux_tree_tapbuf_size2 mux_top_track_304 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[153]}),
		.sram(mux_tree_tapbuf_size2_31_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_31_sram_inv[0:1]),
		.out(chany_top_out[152]));

	mux_tree_tapbuf_size2 mux_top_track_320 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[161]}),
		.sram(mux_tree_tapbuf_size2_32_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_32_sram_inv[0:1]),
		.out(chany_top_out[160]));

	mux_tree_tapbuf_size2 mux_top_track_322 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[162]}),
		.sram(mux_tree_tapbuf_size2_33_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_33_sram_inv[0:1]),
		.out(chany_top_out[161]));

	mux_tree_tapbuf_size2 mux_top_track_338 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[170]}),
		.sram(mux_tree_tapbuf_size2_34_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_34_sram_inv[0:1]),
		.out(chany_top_out[169]));

	mux_tree_tapbuf_size2 mux_top_track_340 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[171]}),
		.sram(mux_tree_tapbuf_size2_35_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_35_sram_inv[0:1]),
		.out(chany_top_out[170]));

	mux_tree_tapbuf_size2 mux_top_track_356 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[179]}),
		.sram(mux_tree_tapbuf_size2_36_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_36_sram_inv[0:1]),
		.out(chany_top_out[178]));

	mux_tree_tapbuf_size2 mux_top_track_358 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[180]}),
		.sram(mux_tree_tapbuf_size2_37_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_37_sram_inv[0:1]),
		.out(chany_top_out[179]));

	mux_tree_tapbuf_size2 mux_top_track_374 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[188]}),
		.sram(mux_tree_tapbuf_size2_38_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_38_sram_inv[0:1]),
		.out(chany_top_out[187]));

	mux_tree_tapbuf_size2 mux_top_track_376 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[189]}),
		.sram(mux_tree_tapbuf_size2_39_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_39_sram_inv[0:1]),
		.out(chany_top_out[188]));

	mux_tree_tapbuf_size2 mux_top_track_392 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[197]}),
		.sram(mux_tree_tapbuf_size2_40_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_40_sram_inv[0:1]),
		.out(chany_top_out[196]));

	mux_tree_tapbuf_size2 mux_top_track_394 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[198]}),
		.sram(mux_tree_tapbuf_size2_41_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_41_sram_inv[0:1]),
		.out(chany_top_out[197]));

	mux_tree_tapbuf_size2 mux_top_track_410 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[206]}),
		.sram(mux_tree_tapbuf_size2_42_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_42_sram_inv[0:1]),
		.out(chany_top_out[205]));

	mux_tree_tapbuf_size2 mux_top_track_412 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[207]}),
		.sram(mux_tree_tapbuf_size2_43_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_43_sram_inv[0:1]),
		.out(chany_top_out[206]));

	mux_tree_tapbuf_size2 mux_top_track_428 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[215]}),
		.sram(mux_tree_tapbuf_size2_44_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_44_sram_inv[0:1]),
		.out(chany_top_out[214]));

	mux_tree_tapbuf_size2 mux_top_track_430 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[216]}),
		.sram(mux_tree_tapbuf_size2_45_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_45_sram_inv[0:1]),
		.out(chany_top_out[215]));

	mux_tree_tapbuf_size2 mux_top_track_446 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[224]}),
		.sram(mux_tree_tapbuf_size2_46_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_46_sram_inv[0:1]),
		.out(chany_top_out[223]));

	mux_tree_tapbuf_size2 mux_top_track_448 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[225]}),
		.sram(mux_tree_tapbuf_size2_47_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_47_sram_inv[0:1]),
		.out(chany_top_out[224]));

	mux_tree_tapbuf_size2 mux_top_track_464 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[233]}),
		.sram(mux_tree_tapbuf_size2_48_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_48_sram_inv[0:1]),
		.out(chany_top_out[232]));

	mux_tree_tapbuf_size2 mux_top_track_466 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[234]}),
		.sram(mux_tree_tapbuf_size2_49_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_49_sram_inv[0:1]),
		.out(chany_top_out[233]));

	mux_tree_tapbuf_size2 mux_top_track_482 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[242]}),
		.sram(mux_tree_tapbuf_size2_50_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_50_sram_inv[0:1]),
		.out(chany_top_out[241]));

	mux_tree_tapbuf_size2 mux_top_track_484 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[243]}),
		.sram(mux_tree_tapbuf_size2_51_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_51_sram_inv[0:1]),
		.out(chany_top_out[242]));

	mux_tree_tapbuf_size2 mux_top_track_500 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[251]}),
		.sram(mux_tree_tapbuf_size2_52_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_52_sram_inv[0:1]),
		.out(chany_top_out[250]));

	mux_tree_tapbuf_size2 mux_top_track_502 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[252]}),
		.sram(mux_tree_tapbuf_size2_53_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_53_sram_inv[0:1]),
		.out(chany_top_out[251]));

	mux_tree_tapbuf_size2 mux_top_track_518 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[260]}),
		.sram(mux_tree_tapbuf_size2_54_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_54_sram_inv[0:1]),
		.out(chany_top_out[259]));

	mux_tree_tapbuf_size2 mux_top_track_520 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[261]}),
		.sram(mux_tree_tapbuf_size2_55_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_55_sram_inv[0:1]),
		.out(chany_top_out[260]));

	mux_tree_tapbuf_size2 mux_top_track_536 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[269]}),
		.sram(mux_tree_tapbuf_size2_56_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_56_sram_inv[0:1]),
		.out(chany_top_out[268]));

	mux_tree_tapbuf_size2 mux_top_track_538 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[270]}),
		.sram(mux_tree_tapbuf_size2_57_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_57_sram_inv[0:1]),
		.out(chany_top_out[269]));

	mux_tree_tapbuf_size2 mux_top_track_554 (
		.in({top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, chanx_right_in[278]}),
		.sram(mux_tree_tapbuf_size2_58_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_58_sram_inv[0:1]),
		.out(chany_top_out[277]));

	mux_tree_tapbuf_size2 mux_top_track_556 (
		.in({top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_, chanx_right_in[279]}),
		.sram(mux_tree_tapbuf_size2_59_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_59_sram_inv[0:1]),
		.out(chany_top_out[278]));

	mux_tree_tapbuf_size2 mux_right_track_32 (
		.in({chany_top_in[15], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_60_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_60_sram_inv[0:1]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size2 mux_right_track_34 (
		.in({chany_top_in[16], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_61_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_61_sram_inv[0:1]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size2 mux_right_track_50 (
		.in({chany_top_in[24], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_62_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_62_sram_inv[0:1]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size2 mux_right_track_52 (
		.in({chany_top_in[25], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_63_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_63_sram_inv[0:1]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size2 mux_right_track_68 (
		.in({chany_top_in[33], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_64_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_64_sram_inv[0:1]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size2 mux_right_track_70 (
		.in({chany_top_in[34], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_65_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_65_sram_inv[0:1]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size2 mux_right_track_86 (
		.in({chany_top_in[42], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_66_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_66_sram_inv[0:1]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size2 mux_right_track_88 (
		.in({chany_top_in[43], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_67_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_67_sram_inv[0:1]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size2 mux_right_track_104 (
		.in({chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_68_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_68_sram_inv[0:1]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size2 mux_right_track_106 (
		.in({chany_top_in[52], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_69_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_69_sram_inv[0:1]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size2 mux_right_track_122 (
		.in({chany_top_in[60], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_70_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_70_sram_inv[0:1]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size2 mux_right_track_124 (
		.in({chany_top_in[61], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_71_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_71_sram_inv[0:1]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size2 mux_right_track_140 (
		.in({chany_top_in[69], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_72_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_72_sram_inv[0:1]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size2 mux_right_track_142 (
		.in({chany_top_in[70], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_73_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_73_sram_inv[0:1]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size2 mux_right_track_158 (
		.in({chany_top_in[78], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_74_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_74_sram_inv[0:1]),
		.out(chanx_right_out[79]));

	mux_tree_tapbuf_size2 mux_right_track_160 (
		.in({chany_top_in[79], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_75_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_75_sram_inv[0:1]),
		.out(chanx_right_out[80]));

	mux_tree_tapbuf_size2 mux_right_track_176 (
		.in({chany_top_in[87], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_76_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_76_sram_inv[0:1]),
		.out(chanx_right_out[88]));

	mux_tree_tapbuf_size2 mux_right_track_178 (
		.in({chany_top_in[88], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_77_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_77_sram_inv[0:1]),
		.out(chanx_right_out[89]));

	mux_tree_tapbuf_size2 mux_right_track_194 (
		.in({chany_top_in[96], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_78_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_78_sram_inv[0:1]),
		.out(chanx_right_out[97]));

	mux_tree_tapbuf_size2 mux_right_track_196 (
		.in({chany_top_in[97], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_79_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_79_sram_inv[0:1]),
		.out(chanx_right_out[98]));

	mux_tree_tapbuf_size2 mux_right_track_212 (
		.in({chany_top_in[105], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_80_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_80_sram_inv[0:1]),
		.out(chanx_right_out[106]));

	mux_tree_tapbuf_size2 mux_right_track_214 (
		.in({chany_top_in[106], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_81_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_81_sram_inv[0:1]),
		.out(chanx_right_out[107]));

	mux_tree_tapbuf_size2 mux_right_track_230 (
		.in({chany_top_in[114], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_82_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_82_sram_inv[0:1]),
		.out(chanx_right_out[115]));

	mux_tree_tapbuf_size2 mux_right_track_232 (
		.in({chany_top_in[115], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_83_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_83_sram_inv[0:1]),
		.out(chanx_right_out[116]));

	mux_tree_tapbuf_size2 mux_right_track_248 (
		.in({chany_top_in[123], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_84_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_84_sram_inv[0:1]),
		.out(chanx_right_out[124]));

	mux_tree_tapbuf_size2 mux_right_track_250 (
		.in({chany_top_in[124], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_85_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_85_sram_inv[0:1]),
		.out(chanx_right_out[125]));

	mux_tree_tapbuf_size2 mux_right_track_266 (
		.in({chany_top_in[132], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_86_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_86_sram_inv[0:1]),
		.out(chanx_right_out[133]));

	mux_tree_tapbuf_size2 mux_right_track_268 (
		.in({chany_top_in[133], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_87_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_87_sram_inv[0:1]),
		.out(chanx_right_out[134]));

	mux_tree_tapbuf_size2 mux_right_track_284 (
		.in({chany_top_in[141], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_88_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_88_sram_inv[0:1]),
		.out(chanx_right_out[142]));

	mux_tree_tapbuf_size2 mux_right_track_286 (
		.in({chany_top_in[142], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_89_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_89_sram_inv[0:1]),
		.out(chanx_right_out[143]));

	mux_tree_tapbuf_size2 mux_right_track_302 (
		.in({chany_top_in[150], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_90_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_90_sram_inv[0:1]),
		.out(chanx_right_out[151]));

	mux_tree_tapbuf_size2 mux_right_track_304 (
		.in({chany_top_in[151], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_91_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_91_sram_inv[0:1]),
		.out(chanx_right_out[152]));

	mux_tree_tapbuf_size2 mux_right_track_320 (
		.in({chany_top_in[159], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_92_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_92_sram_inv[0:1]),
		.out(chanx_right_out[160]));

	mux_tree_tapbuf_size2 mux_right_track_322 (
		.in({chany_top_in[160], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_93_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_93_sram_inv[0:1]),
		.out(chanx_right_out[161]));

	mux_tree_tapbuf_size2 mux_right_track_338 (
		.in({chany_top_in[168], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_94_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_94_sram_inv[0:1]),
		.out(chanx_right_out[169]));

	mux_tree_tapbuf_size2 mux_right_track_340 (
		.in({chany_top_in[169], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_95_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_95_sram_inv[0:1]),
		.out(chanx_right_out[170]));

	mux_tree_tapbuf_size2 mux_right_track_356 (
		.in({chany_top_in[177], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_96_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_96_sram_inv[0:1]),
		.out(chanx_right_out[178]));

	mux_tree_tapbuf_size2 mux_right_track_358 (
		.in({chany_top_in[178], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_97_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_97_sram_inv[0:1]),
		.out(chanx_right_out[179]));

	mux_tree_tapbuf_size2 mux_right_track_374 (
		.in({chany_top_in[186], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_98_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_98_sram_inv[0:1]),
		.out(chanx_right_out[187]));

	mux_tree_tapbuf_size2 mux_right_track_376 (
		.in({chany_top_in[187], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_99_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_99_sram_inv[0:1]),
		.out(chanx_right_out[188]));

	mux_tree_tapbuf_size2 mux_right_track_392 (
		.in({chany_top_in[195], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_100_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_100_sram_inv[0:1]),
		.out(chanx_right_out[196]));

	mux_tree_tapbuf_size2 mux_right_track_394 (
		.in({chany_top_in[196], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_101_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_101_sram_inv[0:1]),
		.out(chanx_right_out[197]));

	mux_tree_tapbuf_size2 mux_right_track_410 (
		.in({chany_top_in[204], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_102_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_102_sram_inv[0:1]),
		.out(chanx_right_out[205]));

	mux_tree_tapbuf_size2 mux_right_track_412 (
		.in({chany_top_in[205], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_103_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_103_sram_inv[0:1]),
		.out(chanx_right_out[206]));

	mux_tree_tapbuf_size2 mux_right_track_428 (
		.in({chany_top_in[213], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_104_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_104_sram_inv[0:1]),
		.out(chanx_right_out[214]));

	mux_tree_tapbuf_size2 mux_right_track_430 (
		.in({chany_top_in[214], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_105_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_105_sram_inv[0:1]),
		.out(chanx_right_out[215]));

	mux_tree_tapbuf_size2 mux_right_track_446 (
		.in({chany_top_in[222], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_106_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_106_sram_inv[0:1]),
		.out(chanx_right_out[223]));

	mux_tree_tapbuf_size2 mux_right_track_448 (
		.in({chany_top_in[223], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_107_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_107_sram_inv[0:1]),
		.out(chanx_right_out[224]));

	mux_tree_tapbuf_size2 mux_right_track_464 (
		.in({chany_top_in[231], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_108_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_108_sram_inv[0:1]),
		.out(chanx_right_out[232]));

	mux_tree_tapbuf_size2 mux_right_track_466 (
		.in({chany_top_in[232], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_109_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_109_sram_inv[0:1]),
		.out(chanx_right_out[233]));

	mux_tree_tapbuf_size2 mux_right_track_482 (
		.in({chany_top_in[240], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_110_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_110_sram_inv[0:1]),
		.out(chanx_right_out[241]));

	mux_tree_tapbuf_size2 mux_right_track_484 (
		.in({chany_top_in[241], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_111_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_111_sram_inv[0:1]),
		.out(chanx_right_out[242]));

	mux_tree_tapbuf_size2 mux_right_track_500 (
		.in({chany_top_in[249], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_112_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_112_sram_inv[0:1]),
		.out(chanx_right_out[250]));

	mux_tree_tapbuf_size2 mux_right_track_502 (
		.in({chany_top_in[250], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_113_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_113_sram_inv[0:1]),
		.out(chanx_right_out[251]));

	mux_tree_tapbuf_size2 mux_right_track_518 (
		.in({chany_top_in[258], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_114_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_114_sram_inv[0:1]),
		.out(chanx_right_out[259]));

	mux_tree_tapbuf_size2 mux_right_track_520 (
		.in({chany_top_in[259], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_115_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_115_sram_inv[0:1]),
		.out(chanx_right_out[260]));

	mux_tree_tapbuf_size2 mux_right_track_536 (
		.in({chany_top_in[267], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_116_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_116_sram_inv[0:1]),
		.out(chanx_right_out[268]));

	mux_tree_tapbuf_size2 mux_right_track_538 (
		.in({chany_top_in[268], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_117_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_117_sram_inv[0:1]),
		.out(chanx_right_out[269]));

	mux_tree_tapbuf_size2 mux_right_track_554 (
		.in({chany_top_in[276], right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_118_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_118_sram_inv[0:1]),
		.out(chanx_right_out[277]));

	mux_tree_tapbuf_size2 mux_right_track_556 (
		.in({chany_top_in[277], right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size2_119_sram[0:1]),
		.sram_inv(mux_tree_tapbuf_size2_119_sram_inv[0:1]),
		.out(chanx_right_out[278]));

	mux_tree_tapbuf_size2_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_0_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_0_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_1_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_1_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_2_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_2_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_3_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_3_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_4_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_4_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_5_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_5_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_6_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_6_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_7_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_7_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_41_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_8_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_8_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_9_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_9_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_10_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_10_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_11_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_11_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_55_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_12_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_12_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_13_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_13_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_14_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_14_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_15_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_15_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_69_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_16_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_16_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_17_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_17_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_18_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_18_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_19_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_19_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_83_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_20_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_20_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_21_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_21_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_22_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_22_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_23_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_23_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_97_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_24_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_24_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_25_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_25_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_26_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_26_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_27_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_27_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_111_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_28_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_28_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_29_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_29_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_30_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_30_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_31_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_31_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_125_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_32_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_32_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_33_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_33_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_132_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_34_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_34_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_35_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_35_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_139_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_36_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_36_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_37_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_37_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_37_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_146_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_38_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_38_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_38_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_39_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_39_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_39_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_153_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_40_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_40_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_394 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_40_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_41_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_41_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_41_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_410 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_160_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_42_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_42_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_412 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_42_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_43_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_43_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_43_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_428 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_167_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_44_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_44_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_430 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_44_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_45_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_45_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_45_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_446 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_174_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_46_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_46_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_46_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_47_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_47_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_47_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_181_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_48_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_48_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_466 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_48_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_49_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_49_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_49_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_482 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_188_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_50_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_50_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_484 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_50_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_51_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_51_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_51_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_500 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_195_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_52_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_52_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_502 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_52_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_53_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_53_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_53_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_518 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_202_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_54_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_54_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_54_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_55_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_55_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_55_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_209_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_56_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_56_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_538 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_56_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_57_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_57_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_57_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_554 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_216_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_58_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_58_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_top_track_556 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_58_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_59_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_59_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_59_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_236_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_60_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_60_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_60_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_61_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_61_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_61_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_243_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_62_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_62_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_62_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_63_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_63_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_63_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_250_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_64_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_64_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_64_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_65_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_65_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_65_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_257_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_66_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_66_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_66_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_67_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_67_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_67_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_264_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_68_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_68_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_68_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_69_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_69_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_69_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_271_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_70_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_70_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_70_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_71_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_71_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_71_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_278_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_72_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_72_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_72_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_73_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_73_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_73_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_158 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_285_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_74_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_74_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_160 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_74_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_75_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_75_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_75_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_176 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_292_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_76_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_76_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_178 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_76_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_77_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_77_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_77_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_194 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_299_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_78_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_78_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_196 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_78_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_79_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_79_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_79_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_212 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_306_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_80_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_80_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_214 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_80_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_81_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_81_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_81_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_230 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_313_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_82_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_82_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_232 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_82_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_83_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_83_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_83_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_248 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_320_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_84_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_84_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_250 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_84_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_85_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_85_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_85_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_266 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_327_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_86_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_86_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_268 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_86_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_87_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_87_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_87_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_284 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_334_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_88_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_88_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_286 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_88_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_89_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_89_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_89_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_302 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_341_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_90_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_90_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_304 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_90_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_91_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_91_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_91_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_320 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_348_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_92_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_92_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_322 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_92_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_93_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_93_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_93_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_338 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_355_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_94_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_94_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_340 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_94_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_95_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_95_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_95_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_356 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_362_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_96_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_96_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_358 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_96_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_97_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_97_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_97_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_374 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_369_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_98_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_98_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_376 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_98_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_99_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_99_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_99_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_392 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_376_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_100_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_100_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_394 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_100_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_101_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_101_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_101_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_410 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_383_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_102_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_102_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_412 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_102_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_103_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_103_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_103_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_428 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_390_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_104_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_104_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_430 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_104_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_105_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_105_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_105_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_446 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_397_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_106_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_106_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_448 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_106_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_107_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_107_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_107_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_464 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_404_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_108_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_108_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_466 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_108_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_109_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_109_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_109_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_482 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_411_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_110_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_110_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_484 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_110_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_111_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_111_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_111_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_500 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_418_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_112_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_112_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_502 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_112_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_113_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_113_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_113_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_518 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_425_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_114_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_114_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_520 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_114_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_115_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_115_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_115_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_536 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_432_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_116_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_116_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_538 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_116_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_117_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_117_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_117_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_554 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size3_mem_439_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_118_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_118_sram_inv[0:1]));

	mux_tree_tapbuf_size2_mem mem_right_track_556 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size2_mem_118_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size2_mem_119_ccff_tail),
		.mem_out(mux_tree_tapbuf_size2_119_sram[0:1]),
		.mem_outb(mux_tree_tapbuf_size2_119_sram_inv[0:1]));

endmodule
// ----- END Verilog module for sb_0__0_ -----

//----- Default net type -----
`default_nettype wire



