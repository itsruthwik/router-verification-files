//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog modules for Unique Switch Blocks[0][1]
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Sat Jun 29 10:24:45 2024
//-------------------------------------------
//----- Default net type -----
`default_nettype none

// ----- Verilog module for sb_0__1_ -----
module sb_0__1_(prog_clk,
                chany_top_in,
                top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_,
                top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_,
                chanx_right_in,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_,
                right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_,
                right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_,
                chany_bottom_in,
                bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_,
                bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_,
                bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_,
                ccff_head,
                chany_top_out,
                chanx_right_out,
                chany_bottom_out,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- INPUT PORTS -----
input [0:72] chany_top_in;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_;
//----- INPUT PORTS -----
input [0:0] top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_;
//----- INPUT PORTS -----
input [0:72] chanx_right_in;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_;
//----- INPUT PORTS -----
input [0:0] right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_;
//----- INPUT PORTS -----
input [0:0] right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_;
//----- INPUT PORTS -----
input [0:72] chany_bottom_in;
//----- INPUT PORTS -----
input [0:0] bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:72] chany_top_out;
//----- OUTPUT PORTS -----
output [0:72] chanx_right_out;
//----- OUTPUT PORTS -----
output [0:72] chany_bottom_out;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN wire-connection ports -----
//----- END wire-connection ports -----


//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:3] mux_tree_tapbuf_size10_0_sram;
wire [0:3] mux_tree_tapbuf_size10_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size10_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size11_0_sram;
wire [0:3] mux_tree_tapbuf_size11_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_10_sram;
wire [0:3] mux_tree_tapbuf_size11_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_1_sram;
wire [0:3] mux_tree_tapbuf_size11_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_2_sram;
wire [0:3] mux_tree_tapbuf_size11_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_3_sram;
wire [0:3] mux_tree_tapbuf_size11_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_4_sram;
wire [0:3] mux_tree_tapbuf_size11_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_5_sram;
wire [0:3] mux_tree_tapbuf_size11_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_6_sram;
wire [0:3] mux_tree_tapbuf_size11_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_7_sram;
wire [0:3] mux_tree_tapbuf_size11_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_8_sram;
wire [0:3] mux_tree_tapbuf_size11_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size11_9_sram;
wire [0:3] mux_tree_tapbuf_size11_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size11_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size11_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size12_0_sram;
wire [0:3] mux_tree_tapbuf_size12_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_10_sram;
wire [0:3] mux_tree_tapbuf_size12_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_11_sram;
wire [0:3] mux_tree_tapbuf_size12_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_12_sram;
wire [0:3] mux_tree_tapbuf_size12_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_13_sram;
wire [0:3] mux_tree_tapbuf_size12_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_14_sram;
wire [0:3] mux_tree_tapbuf_size12_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_15_sram;
wire [0:3] mux_tree_tapbuf_size12_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_16_sram;
wire [0:3] mux_tree_tapbuf_size12_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_17_sram;
wire [0:3] mux_tree_tapbuf_size12_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_18_sram;
wire [0:3] mux_tree_tapbuf_size12_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_19_sram;
wire [0:3] mux_tree_tapbuf_size12_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_1_sram;
wire [0:3] mux_tree_tapbuf_size12_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_20_sram;
wire [0:3] mux_tree_tapbuf_size12_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_21_sram;
wire [0:3] mux_tree_tapbuf_size12_21_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_22_sram;
wire [0:3] mux_tree_tapbuf_size12_22_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_23_sram;
wire [0:3] mux_tree_tapbuf_size12_23_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_24_sram;
wire [0:3] mux_tree_tapbuf_size12_24_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_25_sram;
wire [0:3] mux_tree_tapbuf_size12_25_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_26_sram;
wire [0:3] mux_tree_tapbuf_size12_26_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_27_sram;
wire [0:3] mux_tree_tapbuf_size12_27_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_28_sram;
wire [0:3] mux_tree_tapbuf_size12_28_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_29_sram;
wire [0:3] mux_tree_tapbuf_size12_29_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_2_sram;
wire [0:3] mux_tree_tapbuf_size12_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_30_sram;
wire [0:3] mux_tree_tapbuf_size12_30_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_31_sram;
wire [0:3] mux_tree_tapbuf_size12_31_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_32_sram;
wire [0:3] mux_tree_tapbuf_size12_32_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_33_sram;
wire [0:3] mux_tree_tapbuf_size12_33_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_34_sram;
wire [0:3] mux_tree_tapbuf_size12_34_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_35_sram;
wire [0:3] mux_tree_tapbuf_size12_35_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_36_sram;
wire [0:3] mux_tree_tapbuf_size12_36_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_3_sram;
wire [0:3] mux_tree_tapbuf_size12_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_4_sram;
wire [0:3] mux_tree_tapbuf_size12_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_5_sram;
wire [0:3] mux_tree_tapbuf_size12_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_6_sram;
wire [0:3] mux_tree_tapbuf_size12_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_7_sram;
wire [0:3] mux_tree_tapbuf_size12_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_8_sram;
wire [0:3] mux_tree_tapbuf_size12_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size12_9_sram;
wire [0:3] mux_tree_tapbuf_size12_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size12_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_21_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_22_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_23_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_24_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_25_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_26_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_27_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_28_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_29_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_30_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_31_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_32_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_33_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_34_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_35_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_36_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size12_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size13_0_sram;
wire [0:3] mux_tree_tapbuf_size13_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_10_sram;
wire [0:3] mux_tree_tapbuf_size13_10_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_11_sram;
wire [0:3] mux_tree_tapbuf_size13_11_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_12_sram;
wire [0:3] mux_tree_tapbuf_size13_12_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_13_sram;
wire [0:3] mux_tree_tapbuf_size13_13_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_14_sram;
wire [0:3] mux_tree_tapbuf_size13_14_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_15_sram;
wire [0:3] mux_tree_tapbuf_size13_15_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_16_sram;
wire [0:3] mux_tree_tapbuf_size13_16_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_17_sram;
wire [0:3] mux_tree_tapbuf_size13_17_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_18_sram;
wire [0:3] mux_tree_tapbuf_size13_18_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_19_sram;
wire [0:3] mux_tree_tapbuf_size13_19_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_1_sram;
wire [0:3] mux_tree_tapbuf_size13_1_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_20_sram;
wire [0:3] mux_tree_tapbuf_size13_20_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_2_sram;
wire [0:3] mux_tree_tapbuf_size13_2_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_3_sram;
wire [0:3] mux_tree_tapbuf_size13_3_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_4_sram;
wire [0:3] mux_tree_tapbuf_size13_4_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_5_sram;
wire [0:3] mux_tree_tapbuf_size13_5_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_6_sram;
wire [0:3] mux_tree_tapbuf_size13_6_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_7_sram;
wire [0:3] mux_tree_tapbuf_size13_7_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_8_sram;
wire [0:3] mux_tree_tapbuf_size13_8_sram_inv;
wire [0:3] mux_tree_tapbuf_size13_9_sram;
wire [0:3] mux_tree_tapbuf_size13_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size13_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_11_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_12_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_13_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_14_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_15_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_16_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_17_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_18_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_19_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_20_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size13_mem_9_ccff_tail;
wire [0:3] mux_tree_tapbuf_size14_0_sram;
wire [0:3] mux_tree_tapbuf_size14_0_sram_inv;
wire [0:3] mux_tree_tapbuf_size14_1_sram;
wire [0:3] mux_tree_tapbuf_size14_1_sram_inv;
wire [0:0] mux_tree_tapbuf_size14_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size14_mem_1_ccff_tail;
wire [0:4] mux_tree_tapbuf_size20_0_sram;
wire [0:4] mux_tree_tapbuf_size20_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_1_sram;
wire [0:4] mux_tree_tapbuf_size20_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_2_sram;
wire [0:4] mux_tree_tapbuf_size20_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_3_sram;
wire [0:4] mux_tree_tapbuf_size20_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_4_sram;
wire [0:4] mux_tree_tapbuf_size20_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size20_5_sram;
wire [0:4] mux_tree_tapbuf_size20_5_sram_inv;
wire [0:0] mux_tree_tapbuf_size20_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size20_mem_5_ccff_tail;
wire [0:4] mux_tree_tapbuf_size21_0_sram;
wire [0:4] mux_tree_tapbuf_size21_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_1_sram;
wire [0:4] mux_tree_tapbuf_size21_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_2_sram;
wire [0:4] mux_tree_tapbuf_size21_2_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_3_sram;
wire [0:4] mux_tree_tapbuf_size21_3_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_4_sram;
wire [0:4] mux_tree_tapbuf_size21_4_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_5_sram;
wire [0:4] mux_tree_tapbuf_size21_5_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_6_sram;
wire [0:4] mux_tree_tapbuf_size21_6_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_7_sram;
wire [0:4] mux_tree_tapbuf_size21_7_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_8_sram;
wire [0:4] mux_tree_tapbuf_size21_8_sram_inv;
wire [0:4] mux_tree_tapbuf_size21_9_sram;
wire [0:4] mux_tree_tapbuf_size21_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size21_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size21_mem_9_ccff_tail;
wire [0:4] mux_tree_tapbuf_size22_0_sram;
wire [0:4] mux_tree_tapbuf_size22_0_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_1_sram;
wire [0:4] mux_tree_tapbuf_size22_1_sram_inv;
wire [0:4] mux_tree_tapbuf_size22_2_sram;
wire [0:4] mux_tree_tapbuf_size22_2_sram_inv;
wire [0:0] mux_tree_tapbuf_size22_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size22_mem_2_ccff_tail;
wire [0:2] mux_tree_tapbuf_size5_0_sram;
wire [0:2] mux_tree_tapbuf_size5_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_1_sram;
wire [0:2] mux_tree_tapbuf_size5_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_2_sram;
wire [0:2] mux_tree_tapbuf_size5_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_3_sram;
wire [0:2] mux_tree_tapbuf_size5_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_4_sram;
wire [0:2] mux_tree_tapbuf_size5_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_5_sram;
wire [0:2] mux_tree_tapbuf_size5_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size5_6_sram;
wire [0:2] mux_tree_tapbuf_size5_6_sram_inv;
wire [0:0] mux_tree_tapbuf_size5_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size5_mem_5_ccff_tail;
wire [0:2] mux_tree_tapbuf_size6_0_sram;
wire [0:2] mux_tree_tapbuf_size6_0_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_10_sram;
wire [0:2] mux_tree_tapbuf_size6_10_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_1_sram;
wire [0:2] mux_tree_tapbuf_size6_1_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_2_sram;
wire [0:2] mux_tree_tapbuf_size6_2_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_3_sram;
wire [0:2] mux_tree_tapbuf_size6_3_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_4_sram;
wire [0:2] mux_tree_tapbuf_size6_4_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_5_sram;
wire [0:2] mux_tree_tapbuf_size6_5_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_6_sram;
wire [0:2] mux_tree_tapbuf_size6_6_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_7_sram;
wire [0:2] mux_tree_tapbuf_size6_7_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_8_sram;
wire [0:2] mux_tree_tapbuf_size6_8_sram_inv;
wire [0:2] mux_tree_tapbuf_size6_9_sram;
wire [0:2] mux_tree_tapbuf_size6_9_sram_inv;
wire [0:0] mux_tree_tapbuf_size6_mem_0_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_10_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_1_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_2_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_3_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_4_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_5_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_6_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_7_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_8_ccff_tail;
wire [0:0] mux_tree_tapbuf_size6_mem_9_ccff_tail;
wire [0:2] mux_tree_tapbuf_size7_0_sram;
wire [0:2] mux_tree_tapbuf_size7_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size7_mem_0_ccff_tail;
wire [0:3] mux_tree_tapbuf_size9_0_sram;
wire [0:3] mux_tree_tapbuf_size9_0_sram_inv;
wire [0:0] mux_tree_tapbuf_size9_mem_0_ccff_tail;

// ----- BEGIN Local short connections -----
// ----- Local connection due to Wire 0 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[1] = chany_top_in[0];
// ----- Local connection due to Wire 1 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[2] = chany_top_in[1];
// ----- Local connection due to Wire 2 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[3] = chany_top_in[2];
// ----- Local connection due to Wire 4 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[5] = chany_top_in[4];
// ----- Local connection due to Wire 5 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[6] = chany_top_in[5];
// ----- Local connection due to Wire 6 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[7] = chany_top_in[6];
// ----- Local connection due to Wire 8 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[9] = chany_top_in[8];
// ----- Local connection due to Wire 9 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[10] = chany_top_in[9];
// ----- Local connection due to Wire 10 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[11] = chany_top_in[10];
// ----- Local connection due to Wire 12 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[13] = chany_top_in[12];
// ----- Local connection due to Wire 13 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[14] = chany_top_in[13];
// ----- Local connection due to Wire 14 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[15] = chany_top_in[14];
// ----- Local connection due to Wire 16 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[17] = chany_top_in[16];
// ----- Local connection due to Wire 17 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[18] = chany_top_in[17];
// ----- Local connection due to Wire 18 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[19] = chany_top_in[18];
// ----- Local connection due to Wire 20 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[21] = chany_top_in[20];
// ----- Local connection due to Wire 21 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[22] = chany_top_in[21];
// ----- Local connection due to Wire 22 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[23] = chany_top_in[22];
// ----- Local connection due to Wire 24 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[25] = chany_top_in[24];
// ----- Local connection due to Wire 25 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[26] = chany_top_in[25];
// ----- Local connection due to Wire 26 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[27] = chany_top_in[26];
// ----- Local connection due to Wire 28 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[29] = chany_top_in[28];
// ----- Local connection due to Wire 29 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[30] = chany_top_in[29];
// ----- Local connection due to Wire 30 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[31] = chany_top_in[30];
// ----- Local connection due to Wire 32 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[33] = chany_top_in[32];
// ----- Local connection due to Wire 33 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[34] = chany_top_in[33];
// ----- Local connection due to Wire 34 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[35] = chany_top_in[34];
// ----- Local connection due to Wire 36 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[37] = chany_top_in[36];
// ----- Local connection due to Wire 37 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[38] = chany_top_in[37];
// ----- Local connection due to Wire 38 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[39] = chany_top_in[38];
// ----- Local connection due to Wire 40 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[41] = chany_top_in[40];
// ----- Local connection due to Wire 41 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[42] = chany_top_in[41];
// ----- Local connection due to Wire 42 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[43] = chany_top_in[42];
// ----- Local connection due to Wire 44 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[45] = chany_top_in[44];
// ----- Local connection due to Wire 45 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[46] = chany_top_in[45];
// ----- Local connection due to Wire 46 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[47] = chany_top_in[46];
// ----- Local connection due to Wire 48 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[49] = chany_top_in[48];
// ----- Local connection due to Wire 49 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[50] = chany_top_in[49];
// ----- Local connection due to Wire 50 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[51] = chany_top_in[50];
// ----- Local connection due to Wire 52 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[53] = chany_top_in[52];
// ----- Local connection due to Wire 53 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[54] = chany_top_in[53];
// ----- Local connection due to Wire 54 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[55] = chany_top_in[54];
// ----- Local connection due to Wire 56 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[57] = chany_top_in[56];
// ----- Local connection due to Wire 57 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[58] = chany_top_in[57];
// ----- Local connection due to Wire 58 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[59] = chany_top_in[58];
// ----- Local connection due to Wire 60 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[61] = chany_top_in[60];
// ----- Local connection due to Wire 61 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[62] = chany_top_in[61];
// ----- Local connection due to Wire 62 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[63] = chany_top_in[62];
// ----- Local connection due to Wire 64 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[65] = chany_top_in[64];
// ----- Local connection due to Wire 65 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[66] = chany_top_in[65];
// ----- Local connection due to Wire 66 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[67] = chany_top_in[66];
// ----- Local connection due to Wire 68 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[69] = chany_top_in[68];
// ----- Local connection due to Wire 69 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[70] = chany_top_in[69];
// ----- Local connection due to Wire 70 -----
// ----- Net source id 0 -----
// ----- Net sink id 1 -----
	assign chany_bottom_out[71] = chany_top_in[70];
// ----- Local connection due to Wire 331 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[1] = chany_bottom_in[0];
// ----- Local connection due to Wire 332 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[2] = chany_bottom_in[1];
// ----- Local connection due to Wire 333 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[3] = chany_bottom_in[2];
// ----- Local connection due to Wire 335 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[5] = chany_bottom_in[4];
// ----- Local connection due to Wire 336 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[6] = chany_bottom_in[5];
// ----- Local connection due to Wire 337 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[7] = chany_bottom_in[6];
// ----- Local connection due to Wire 339 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[9] = chany_bottom_in[8];
// ----- Local connection due to Wire 340 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[10] = chany_bottom_in[9];
// ----- Local connection due to Wire 341 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[11] = chany_bottom_in[10];
// ----- Local connection due to Wire 343 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[13] = chany_bottom_in[12];
// ----- Local connection due to Wire 344 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[14] = chany_bottom_in[13];
// ----- Local connection due to Wire 345 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[15] = chany_bottom_in[14];
// ----- Local connection due to Wire 347 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[17] = chany_bottom_in[16];
// ----- Local connection due to Wire 348 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[18] = chany_bottom_in[17];
// ----- Local connection due to Wire 349 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[19] = chany_bottom_in[18];
// ----- Local connection due to Wire 351 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[21] = chany_bottom_in[20];
// ----- Local connection due to Wire 352 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[22] = chany_bottom_in[21];
// ----- Local connection due to Wire 353 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[23] = chany_bottom_in[22];
// ----- Local connection due to Wire 355 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[25] = chany_bottom_in[24];
// ----- Local connection due to Wire 356 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[26] = chany_bottom_in[25];
// ----- Local connection due to Wire 357 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[27] = chany_bottom_in[26];
// ----- Local connection due to Wire 359 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[29] = chany_bottom_in[28];
// ----- Local connection due to Wire 360 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[30] = chany_bottom_in[29];
// ----- Local connection due to Wire 361 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[31] = chany_bottom_in[30];
// ----- Local connection due to Wire 363 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[33] = chany_bottom_in[32];
// ----- Local connection due to Wire 364 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[34] = chany_bottom_in[33];
// ----- Local connection due to Wire 365 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[35] = chany_bottom_in[34];
// ----- Local connection due to Wire 367 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[37] = chany_bottom_in[36];
// ----- Local connection due to Wire 368 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[38] = chany_bottom_in[37];
// ----- Local connection due to Wire 369 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[39] = chany_bottom_in[38];
// ----- Local connection due to Wire 371 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[41] = chany_bottom_in[40];
// ----- Local connection due to Wire 372 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[42] = chany_bottom_in[41];
// ----- Local connection due to Wire 373 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[43] = chany_bottom_in[42];
// ----- Local connection due to Wire 375 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[45] = chany_bottom_in[44];
// ----- Local connection due to Wire 376 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[46] = chany_bottom_in[45];
// ----- Local connection due to Wire 377 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[47] = chany_bottom_in[46];
// ----- Local connection due to Wire 379 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[49] = chany_bottom_in[48];
// ----- Local connection due to Wire 380 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[50] = chany_bottom_in[49];
// ----- Local connection due to Wire 381 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[51] = chany_bottom_in[50];
// ----- Local connection due to Wire 383 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[53] = chany_bottom_in[52];
// ----- Local connection due to Wire 384 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[54] = chany_bottom_in[53];
// ----- Local connection due to Wire 385 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[55] = chany_bottom_in[54];
// ----- Local connection due to Wire 387 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[57] = chany_bottom_in[56];
// ----- Local connection due to Wire 388 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[58] = chany_bottom_in[57];
// ----- Local connection due to Wire 389 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[59] = chany_bottom_in[58];
// ----- Local connection due to Wire 391 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[61] = chany_bottom_in[60];
// ----- Local connection due to Wire 392 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[62] = chany_bottom_in[61];
// ----- Local connection due to Wire 393 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[63] = chany_bottom_in[62];
// ----- Local connection due to Wire 395 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[65] = chany_bottom_in[64];
// ----- Local connection due to Wire 396 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[66] = chany_bottom_in[65];
// ----- Local connection due to Wire 397 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[67] = chany_bottom_in[66];
// ----- Local connection due to Wire 399 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[69] = chany_bottom_in[68];
// ----- Local connection due to Wire 400 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[70] = chany_bottom_in[69];
// ----- Local connection due to Wire 401 -----
// ----- Net source id 0 -----
// ----- Net sink id 0 -----
	assign chany_top_out[71] = chany_bottom_in[70];
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	mux_tree_tapbuf_size22 mux_top_track_0 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[1], chanx_right_in[20], chanx_right_in[39], chanx_right_in[58]}),
		.sram(mux_tree_tapbuf_size22_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_0_sram_inv[0:4]),
		.out(chany_top_out[0]));

	mux_tree_tapbuf_size22 mux_top_track_48 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[7], chanx_right_in[26], chanx_right_in[45], chanx_right_in[64]}),
		.sram(mux_tree_tapbuf_size22_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_1_sram_inv[0:4]),
		.out(chany_top_out[24]));

	mux_tree_tapbuf_size22 mux_top_track_144 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[0], chanx_right_in[19], chanx_right_in[38], chanx_right_in[57]}),
		.sram(mux_tree_tapbuf_size22_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size22_2_sram_inv[0:4]),
		.out(chany_top_out[72]));

	mux_tree_tapbuf_size22_mem mem_top_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(ccff_head),
		.ccff_tail(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_0_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_top_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_1_sram_inv[0:4]));

	mux_tree_tapbuf_size22_mem mem_top_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size22_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size22_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size22_2_sram_inv[0:4]));

	mux_tree_tapbuf_size21 mux_top_track_8 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, chanx_right_in[2], chanx_right_in[21], chanx_right_in[40], chanx_right_in[59]}),
		.sram(mux_tree_tapbuf_size21_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_0_sram_inv[0:4]),
		.out(chany_top_out[4]));

	mux_tree_tapbuf_size21 mux_top_track_32 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[5], chanx_right_in[24], chanx_right_in[43], chanx_right_in[62]}),
		.sram(mux_tree_tapbuf_size21_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_1_sram_inv[0:4]),
		.out(chany_top_out[16]));

	mux_tree_tapbuf_size21 mux_top_track_40 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[6], chanx_right_in[25], chanx_right_in[44], chanx_right_in[63]}),
		.sram(mux_tree_tapbuf_size21_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_2_sram_inv[0:4]),
		.out(chany_top_out[20]));

	mux_tree_tapbuf_size21 mux_top_track_56 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, chanx_right_in[8], chanx_right_in[27], chanx_right_in[46], chanx_right_in[65]}),
		.sram(mux_tree_tapbuf_size21_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_3_sram_inv[0:4]),
		.out(chany_top_out[28]));

	mux_tree_tapbuf_size21 mux_top_track_64 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[9], chanx_right_in[28], chanx_right_in[47], chanx_right_in[66]}),
		.sram(mux_tree_tapbuf_size21_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_4_sram_inv[0:4]),
		.out(chany_top_out[32]));

	mux_tree_tapbuf_size21 mux_top_track_72 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_121_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_157_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_197_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_233_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_273_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_309_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_9_, chanx_right_in[10], chanx_right_in[29], chanx_right_in[48], chanx_right_in[67]}),
		.sram(mux_tree_tapbuf_size21_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_5_sram_inv[0:4]),
		.out(chany_top_out[36]));

	mux_tree_tapbuf_size21 mux_top_track_80 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_125_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_161_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_201_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_237_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_277_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_313_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[11], chanx_right_in[30], chanx_right_in[49], chanx_right_in[68]}),
		.sram(mux_tree_tapbuf_size21_6_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_6_sram_inv[0:4]),
		.out(chany_top_out[40]));

	mux_tree_tapbuf_size21 mux_top_track_96 (
		.in({top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_45_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_69_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[13], chanx_right_in[32], chanx_right_in[51], chanx_right_in[70]}),
		.sram(mux_tree_tapbuf_size21_7_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_7_sram_inv[0:4]),
		.out(chany_top_out[48]));

	mux_tree_tapbuf_size21 mux_top_track_104 (
		.in({top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_21_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_49_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_73_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_97_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, chanx_right_in[14], chanx_right_in[33], chanx_right_in[52], chanx_right_in[71]}),
		.sram(mux_tree_tapbuf_size21_8_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_8_sram_inv[0:4]),
		.out(chany_top_out[52]));

	mux_tree_tapbuf_size21 mux_top_track_112 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_25_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_77_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_101_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_141_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_177_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_217_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_253_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_293_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_329_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, chanx_right_in[15], chanx_right_in[34], chanx_right_in[53], chanx_right_in[72]}),
		.sram(mux_tree_tapbuf_size21_9_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size21_9_sram_inv[0:4]),
		.out(chany_top_out[56]));

	mux_tree_tapbuf_size21_mem mem_top_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_0_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_1_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_2_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_3_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_4_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_5_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_6_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_6_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_7_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_7_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_8_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_8_sram_inv[0:4]));

	mux_tree_tapbuf_size21_mem mem_top_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size21_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size21_9_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size21_9_sram_inv[0:4]));

	mux_tree_tapbuf_size20 mux_top_track_16 (
		.in({top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_53_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[3], chanx_right_in[22], chanx_right_in[41], chanx_right_in[60]}),
		.sram(mux_tree_tapbuf_size20_0_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_0_sram_inv[0:4]),
		.out(chany_top_out[8]));

	mux_tree_tapbuf_size20 mux_top_track_24 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_133_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_137_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_173_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_209_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_213_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_249_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_285_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_289_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_325_, chanx_right_in[4], chanx_right_in[23], chanx_right_in[42], chanx_right_in[61]}),
		.sram(mux_tree_tapbuf_size20_1_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_1_sram_inv[0:4]),
		.out(chany_top_out[12]));

	mux_tree_tapbuf_size20 mux_top_track_88 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_17_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_93_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_129_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_165_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_169_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_205_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_241_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_245_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_281_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_317_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_321_, chanx_right_in[12], chanx_right_in[31], chanx_right_in[50], chanx_right_in[69]}),
		.sram(mux_tree_tapbuf_size20_2_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_2_sram_inv[0:4]),
		.out(chany_top_out[44]));

	mux_tree_tapbuf_size20 mux_top_track_120 (
		.in({top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_5_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_29_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_57_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_81_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_105_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_145_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_181_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_221_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_257_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_297_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_333_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, chanx_right_in[16], chanx_right_in[35], chanx_right_in[54]}),
		.sram(mux_tree_tapbuf_size20_3_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_3_sram_inv[0:4]),
		.out(chany_top_out[60]));

	mux_tree_tapbuf_size20 mux_top_track_128 (
		.in({top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_9_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_33_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_61_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_85_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_109_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_149_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_185_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_225_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_261_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_301_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_337_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, chanx_right_in[17], chanx_right_in[36], chanx_right_in[55]}),
		.sram(mux_tree_tapbuf_size20_4_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_4_sram_inv[0:4]),
		.out(chany_top_out[64]));

	mux_tree_tapbuf_size20 mux_top_track_136 (
		.in({top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_13_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_37_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_41_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_65_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_89_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_113_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_117_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_153_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_189_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_193_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_229_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_265_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_269_, top_right_grid_left_width_0_height_0_subtile_0__pin_channel_out_op_305_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_1_, top_right_grid_left_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_5_, chanx_right_in[18], chanx_right_in[37], chanx_right_in[56]}),
		.sram(mux_tree_tapbuf_size20_5_sram[0:4]),
		.sram_inv(mux_tree_tapbuf_size20_5_sram_inv[0:4]),
		.out(chany_top_out[68]));

	mux_tree_tapbuf_size20_mem mem_top_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_0_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_0_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_top_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_1_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_1_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_top_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_2_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_2_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_top_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size21_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_3_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_3_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_top_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_4_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_4_sram_inv[0:4]));

	mux_tree_tapbuf_size20_mem mem_top_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size20_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size20_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size20_5_sram[0:4]),
		.mem_outb(mux_tree_tapbuf_size20_5_sram_inv[0:4]));

	mux_tree_tapbuf_size11 mux_right_track_0 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size11_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_0_sram_inv[0:3]),
		.out(chanx_right_out[0]));

	mux_tree_tapbuf_size11 mux_right_track_32 (
		.in({chany_top_in[20], chany_top_in[63], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size11_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_1_sram_inv[0:3]),
		.out(chanx_right_out[16]));

	mux_tree_tapbuf_size11 mux_right_track_34 (
		.in({chany_top_in[21], chany_top_in[67], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size11_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_2_sram_inv[0:3]),
		.out(chanx_right_out[17]));

	mux_tree_tapbuf_size11 mux_right_track_44 (
		.in({chany_top_in[28], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[65]}),
		.sram(mux_tree_tapbuf_size11_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_3_sram_inv[0:3]),
		.out(chanx_right_out[22]));

	mux_tree_tapbuf_size11 mux_right_track_52 (
		.in({chany_top_in[33], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[60]}),
		.sram(mux_tree_tapbuf_size11_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_4_sram_inv[0:3]),
		.out(chanx_right_out[26]));

	mux_tree_tapbuf_size11 mux_right_track_64 (
		.in({chany_top_in[41], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[52]}),
		.sram(mux_tree_tapbuf_size11_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_5_sram_inv[0:3]),
		.out(chanx_right_out[32]));

	mux_tree_tapbuf_size11 mux_right_track_70 (
		.in({chany_top_in[45], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[48]}),
		.sram(mux_tree_tapbuf_size11_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_6_sram_inv[0:3]),
		.out(chanx_right_out[35]));

	mux_tree_tapbuf_size11 mux_right_track_84 (
		.in({chany_top_in[54], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[38]}),
		.sram(mux_tree_tapbuf_size11_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_7_sram_inv[0:3]),
		.out(chanx_right_out[42]));

	mux_tree_tapbuf_size11 mux_right_track_88 (
		.in({chany_top_in[57], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[36]}),
		.sram(mux_tree_tapbuf_size11_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_8_sram_inv[0:3]),
		.out(chanx_right_out[44]));

	mux_tree_tapbuf_size11 mux_right_track_104 (
		.in({chany_top_in[68], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[25]}),
		.sram(mux_tree_tapbuf_size11_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_9_sram_inv[0:3]),
		.out(chanx_right_out[52]));

	mux_tree_tapbuf_size11 mux_right_track_142 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[0], chany_bottom_in[3]}),
		.sram(mux_tree_tapbuf_size11_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size11_10_sram_inv[0:3]),
		.out(chanx_right_out[71]));

	mux_tree_tapbuf_size11_mem mem_right_track_0 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size22_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_0_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_32 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_1_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_34 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_2_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_44 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_3_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_52 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_4_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_64 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_5_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_70 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_6_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_84 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_7_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_88 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_8_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_104 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_9_sram_inv[0:3]));

	mux_tree_tapbuf_size11_mem mem_right_track_142 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size11_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size11_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13 mux_right_track_2 (
		.in({chany_top_in[0], chany_top_in[3], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size13_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_0_sram_inv[0:3]),
		.out(chanx_right_out[1]));

	mux_tree_tapbuf_size13 mux_right_track_6 (
		.in({chany_top_in[2], chany_top_in[11], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_}),
		.sram(mux_tree_tapbuf_size13_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_1_sram_inv[0:3]),
		.out(chanx_right_out[3]));

	mux_tree_tapbuf_size13 mux_right_track_8 (
		.in({chany_top_in[4], chany_top_in[15], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_}),
		.sram(mux_tree_tapbuf_size13_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_2_sram_inv[0:3]),
		.out(chanx_right_out[4]));

	mux_tree_tapbuf_size13 mux_right_track_10 (
		.in({chany_top_in[5], chany_top_in[19], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_}),
		.sram(mux_tree_tapbuf_size13_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_3_sram_inv[0:3]),
		.out(chanx_right_out[5]));

	mux_tree_tapbuf_size13 mux_right_track_12 (
		.in({chany_top_in[6], chany_top_in[23], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size13_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_4_sram_inv[0:3]),
		.out(chanx_right_out[6]));

	mux_tree_tapbuf_size13 mux_right_track_20 (
		.in({chany_top_in[12], chany_top_in[39], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_5_sram_inv[0:3]),
		.out(chanx_right_out[10]));

	mux_tree_tapbuf_size13 mux_right_track_24 (
		.in({chany_top_in[14], chany_top_in[47], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size13_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_6_sram_inv[0:3]),
		.out(chanx_right_out[12]));

	mux_tree_tapbuf_size13 mux_right_track_26 (
		.in({chany_top_in[16], chany_top_in[51], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_}),
		.sram(mux_tree_tapbuf_size13_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_7_sram_inv[0:3]),
		.out(chanx_right_out[13]));

	mux_tree_tapbuf_size13 mux_right_track_28 (
		.in({chany_top_in[17], chany_top_in[55], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size13_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_8_sram_inv[0:3]),
		.out(chanx_right_out[14]));

	mux_tree_tapbuf_size13 mux_right_track_30 (
		.in({chany_top_in[18], chany_top_in[59], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size13_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_9_sram_inv[0:3]),
		.out(chanx_right_out[15]));

	mux_tree_tapbuf_size13 mux_right_track_36 (
		.in({chany_top_in[22], chany_top_in[71], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[70]}),
		.sram(mux_tree_tapbuf_size13_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_10_sram_inv[0:3]),
		.out(chanx_right_out[18]));

	mux_tree_tapbuf_size13 mux_right_track_38 (
		.in({chany_top_in[24], chany_top_in[72], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[69]}),
		.sram(mux_tree_tapbuf_size13_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_11_sram_inv[0:3]),
		.out(chanx_right_out[19]));

	mux_tree_tapbuf_size13 mux_right_track_42 (
		.in({chany_top_in[26], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[66]}),
		.sram(mux_tree_tapbuf_size13_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_12_sram_inv[0:3]),
		.out(chanx_right_out[21]));

	mux_tree_tapbuf_size13 mux_right_track_46 (
		.in({chany_top_in[29], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[64]}),
		.sram(mux_tree_tapbuf_size13_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_13_sram_inv[0:3]),
		.out(chanx_right_out[23]));

	mux_tree_tapbuf_size13 mux_right_track_48 (
		.in({chany_top_in[30], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[62]}),
		.sram(mux_tree_tapbuf_size13_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_14_sram_inv[0:3]),
		.out(chanx_right_out[24]));

	mux_tree_tapbuf_size13 mux_right_track_60 (
		.in({chany_top_in[38], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[54]}),
		.sram(mux_tree_tapbuf_size13_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_15_sram_inv[0:3]),
		.out(chanx_right_out[30]));

	mux_tree_tapbuf_size13 mux_right_track_78 (
		.in({chany_top_in[50], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[42]}),
		.sram(mux_tree_tapbuf_size13_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_16_sram_inv[0:3]),
		.out(chanx_right_out[39]));

	mux_tree_tapbuf_size13 mux_right_track_96 (
		.in({chany_top_in[62], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[30]}),
		.sram(mux_tree_tapbuf_size13_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_17_sram_inv[0:3]),
		.out(chanx_right_out[48]));

	mux_tree_tapbuf_size13 mux_right_track_108 (
		.in({chany_top_in[70], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[22], chany_bottom_in[71]}),
		.sram(mux_tree_tapbuf_size13_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_18_sram_inv[0:3]),
		.out(chanx_right_out[54]));

	mux_tree_tapbuf_size13 mux_right_track_114 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[18], chany_bottom_in[59]}),
		.sram(mux_tree_tapbuf_size13_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_19_sram_inv[0:3]),
		.out(chanx_right_out[57]));

	mux_tree_tapbuf_size13 mux_right_track_132 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, chany_bottom_in[6], chany_bottom_in[23]}),
		.sram(mux_tree_tapbuf_size13_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size13_20_sram_inv[0:3]),
		.out(chanx_right_out[66]));

	mux_tree_tapbuf_size13_mem mem_right_track_2 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_0_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_6 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_1_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_8 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_2_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_10 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_3_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_12 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_4_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_20 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_5_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_24 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size14_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_6_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_26 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_7_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_28 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_8_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_30 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_9_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_36 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_10_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_38 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_11_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_42 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_12_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_46 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_13_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_48 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_14_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_60 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_15_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_78 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_16_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_96 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_17_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_108 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_18_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_114 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_19_sram_inv[0:3]));

	mux_tree_tapbuf_size13_mem mem_right_track_132 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size13_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size13_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size13_20_sram_inv[0:3]));

	mux_tree_tapbuf_size14 mux_right_track_4 (
		.in({chany_top_in[1], chany_top_in[7], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_12_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_}),
		.sram(mux_tree_tapbuf_size14_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_0_sram_inv[0:3]),
		.out(chanx_right_out[2]));

	mux_tree_tapbuf_size14 mux_right_track_22 (
		.in({chany_top_in[13], chany_top_in[43], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_48_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_}),
		.sram(mux_tree_tapbuf_size14_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size14_1_sram_inv[0:3]),
		.out(chanx_right_out[11]));

	mux_tree_tapbuf_size14_mem mem_right_track_4 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_0_sram_inv[0:3]));

	mux_tree_tapbuf_size14_mem mem_right_track_22 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size14_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size14_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size14_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12 mux_right_track_14 (
		.in({chany_top_in[8], chany_top_in[27], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_}),
		.sram(mux_tree_tapbuf_size12_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_0_sram_inv[0:3]),
		.out(chanx_right_out[7]));

	mux_tree_tapbuf_size12 mux_right_track_16 (
		.in({chany_top_in[9], chany_top_in[31], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_}),
		.sram(mux_tree_tapbuf_size12_1_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_1_sram_inv[0:3]),
		.out(chanx_right_out[8]));

	mux_tree_tapbuf_size12 mux_right_track_18 (
		.in({chany_top_in[10], chany_top_in[35], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_}),
		.sram(mux_tree_tapbuf_size12_2_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_2_sram_inv[0:3]),
		.out(chanx_right_out[9]));

	mux_tree_tapbuf_size12 mux_right_track_40 (
		.in({chany_top_in[25], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_84_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[68]}),
		.sram(mux_tree_tapbuf_size12_3_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_3_sram_inv[0:3]),
		.out(chanx_right_out[20]));

	mux_tree_tapbuf_size12 mux_right_track_50 (
		.in({chany_top_in[32], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[61]}),
		.sram(mux_tree_tapbuf_size12_4_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_4_sram_inv[0:3]),
		.out(chanx_right_out[25]));

	mux_tree_tapbuf_size12 mux_right_track_54 (
		.in({chany_top_in[34], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[58]}),
		.sram(mux_tree_tapbuf_size12_5_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_5_sram_inv[0:3]),
		.out(chanx_right_out[27]));

	mux_tree_tapbuf_size12 mux_right_track_56 (
		.in({chany_top_in[36], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[57]}),
		.sram(mux_tree_tapbuf_size12_6_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_6_sram_inv[0:3]),
		.out(chanx_right_out[28]));

	mux_tree_tapbuf_size12 mux_right_track_58 (
		.in({chany_top_in[37], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[56]}),
		.sram(mux_tree_tapbuf_size12_7_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_7_sram_inv[0:3]),
		.out(chanx_right_out[29]));

	mux_tree_tapbuf_size12 mux_right_track_62 (
		.in({chany_top_in[40], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[53]}),
		.sram(mux_tree_tapbuf_size12_8_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_8_sram_inv[0:3]),
		.out(chanx_right_out[31]));

	mux_tree_tapbuf_size12 mux_right_track_66 (
		.in({chany_top_in[42], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[50]}),
		.sram(mux_tree_tapbuf_size12_9_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_9_sram_inv[0:3]),
		.out(chanx_right_out[33]));

	mux_tree_tapbuf_size12 mux_right_track_68 (
		.in({chany_top_in[44], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[49]}),
		.sram(mux_tree_tapbuf_size12_10_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_10_sram_inv[0:3]),
		.out(chanx_right_out[34]));

	mux_tree_tapbuf_size12 mux_right_track_72 (
		.in({chany_top_in[46], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[46]}),
		.sram(mux_tree_tapbuf_size12_11_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_11_sram_inv[0:3]),
		.out(chanx_right_out[36]));

	mux_tree_tapbuf_size12 mux_right_track_74 (
		.in({chany_top_in[48], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[45]}),
		.sram(mux_tree_tapbuf_size12_12_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_12_sram_inv[0:3]),
		.out(chanx_right_out[37]));

	mux_tree_tapbuf_size12 mux_right_track_76 (
		.in({chany_top_in[49], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[44]}),
		.sram(mux_tree_tapbuf_size12_13_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_13_sram_inv[0:3]),
		.out(chanx_right_out[38]));

	mux_tree_tapbuf_size12 mux_right_track_80 (
		.in({chany_top_in[52], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[41]}),
		.sram(mux_tree_tapbuf_size12_14_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_14_sram_inv[0:3]),
		.out(chanx_right_out[40]));

	mux_tree_tapbuf_size12 mux_right_track_82 (
		.in({chany_top_in[53], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[40]}),
		.sram(mux_tree_tapbuf_size12_15_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_15_sram_inv[0:3]),
		.out(chanx_right_out[41]));

	mux_tree_tapbuf_size12 mux_right_track_86 (
		.in({chany_top_in[56], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[37]}),
		.sram(mux_tree_tapbuf_size12_16_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_16_sram_inv[0:3]),
		.out(chanx_right_out[43]));

	mux_tree_tapbuf_size12 mux_right_track_90 (
		.in({chany_top_in[58], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[34]}),
		.sram(mux_tree_tapbuf_size12_17_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_17_sram_inv[0:3]),
		.out(chanx_right_out[45]));

	mux_tree_tapbuf_size12 mux_right_track_92 (
		.in({chany_top_in[60], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[33]}),
		.sram(mux_tree_tapbuf_size12_18_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_18_sram_inv[0:3]),
		.out(chanx_right_out[46]));

	mux_tree_tapbuf_size12 mux_right_track_94 (
		.in({chany_top_in[61], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[32]}),
		.sram(mux_tree_tapbuf_size12_19_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_19_sram_inv[0:3]),
		.out(chanx_right_out[47]));

	mux_tree_tapbuf_size12 mux_right_track_98 (
		.in({chany_top_in[64], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[29]}),
		.sram(mux_tree_tapbuf_size12_20_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_20_sram_inv[0:3]),
		.out(chanx_right_out[49]));

	mux_tree_tapbuf_size12 mux_right_track_100 (
		.in({chany_top_in[65], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[28]}),
		.sram(mux_tree_tapbuf_size12_21_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_21_sram_inv[0:3]),
		.out(chanx_right_out[50]));

	mux_tree_tapbuf_size12 mux_right_track_102 (
		.in({chany_top_in[66], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[26]}),
		.sram(mux_tree_tapbuf_size12_22_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_22_sram_inv[0:3]),
		.out(chanx_right_out[51]));

	mux_tree_tapbuf_size12 mux_right_track_106 (
		.in({chany_top_in[69], right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[24], chany_bottom_in[72]}),
		.sram(mux_tree_tapbuf_size12_23_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_23_sram_inv[0:3]),
		.out(chanx_right_out[53]));

	mux_tree_tapbuf_size12 mux_right_track_110 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[21], chany_bottom_in[67]}),
		.sram(mux_tree_tapbuf_size12_24_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_24_sram_inv[0:3]),
		.out(chanx_right_out[55]));

	mux_tree_tapbuf_size12 mux_right_track_112 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_104_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_144_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_184_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_224_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_316_, chany_bottom_in[20], chany_bottom_in[63]}),
		.sram(mux_tree_tapbuf_size12_25_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_25_sram_inv[0:3]),
		.out(chanx_right_out[56]));

	mux_tree_tapbuf_size12 mux_right_track_116 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[17], chany_bottom_in[55]}),
		.sram(mux_tree_tapbuf_size12_26_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_26_sram_inv[0:3]),
		.out(chanx_right_out[58]));

	mux_tree_tapbuf_size12 mux_right_track_118 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[16], chany_bottom_in[51]}),
		.sram(mux_tree_tapbuf_size12_27_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_27_sram_inv[0:3]),
		.out(chanx_right_out[59]));

	mux_tree_tapbuf_size12 mux_right_track_120 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[14], chany_bottom_in[47]}),
		.sram(mux_tree_tapbuf_size12_28_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_28_sram_inv[0:3]),
		.out(chanx_right_out[60]));

	mux_tree_tapbuf_size12 mux_right_track_122 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_124_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_164_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_204_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_244_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_296_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_336_, chany_bottom_in[13], chany_bottom_in[43]}),
		.sram(mux_tree_tapbuf_size12_29_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_29_sram_inv[0:3]),
		.out(chanx_right_out[61]));

	mux_tree_tapbuf_size12 mux_right_track_126 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_132_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_172_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_212_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_252_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_264_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_304_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_4_, chany_bottom_in[10], chany_bottom_in[35]}),
		.sram(mux_tree_tapbuf_size12_30_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_30_sram_inv[0:3]),
		.out(chanx_right_out[63]));

	mux_tree_tapbuf_size12 mux_right_track_128 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_4_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_40_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_76_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_136_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_176_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_216_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_256_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_308_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_flow_ctrl_out_ip_8_, chany_bottom_in[9], chany_bottom_in[31]}),
		.sram(mux_tree_tapbuf_size12_31_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_31_sram_inv[0:3]),
		.out(chanx_right_out[64]));

	mux_tree_tapbuf_size12 mux_right_track_130 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_8_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_44_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_80_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_140_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_180_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_220_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_312_, right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_, chany_bottom_in[8], chany_bottom_in[27]}),
		.sram(mux_tree_tapbuf_size12_32_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_32_sram_inv[0:3]),
		.out(chanx_right_out[65]));

	mux_tree_tapbuf_size12 mux_right_track_134 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_16_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_52_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_88_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_108_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_148_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_188_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_228_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_268_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_320_, chany_bottom_in[5], chany_bottom_in[19]}),
		.sram(mux_tree_tapbuf_size12_33_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_33_sram_inv[0:3]),
		.out(chanx_right_out[67]));

	mux_tree_tapbuf_size12 mux_right_track_136 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_20_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_56_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_92_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_112_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_152_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_192_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_232_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_272_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_284_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_324_, chany_bottom_in[4], chany_bottom_in[15]}),
		.sram(mux_tree_tapbuf_size12_34_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_34_sram_inv[0:3]),
		.out(chanx_right_out[68]));

	mux_tree_tapbuf_size12 mux_right_track_138 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_24_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_60_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_96_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_116_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_156_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_196_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_236_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_276_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_328_, chany_bottom_in[2], chany_bottom_in[11]}),
		.sram(mux_tree_tapbuf_size12_35_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_35_sram_inv[0:3]),
		.out(chanx_right_out[69]));

	mux_tree_tapbuf_size12 mux_right_track_140 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_28_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_64_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_100_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_120_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_160_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_200_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_240_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_280_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_292_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_332_, chany_bottom_in[1], chany_bottom_in[7]}),
		.sram(mux_tree_tapbuf_size12_36_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size12_36_sram_inv[0:3]),
		.out(chanx_right_out[70]));

	mux_tree_tapbuf_size12_mem mem_right_track_14 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_0_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_16 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_1_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_1_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_18 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_2_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_2_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_40 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_3_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_3_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_50 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_4_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_4_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_54 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_5_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_5_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_56 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_6_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_6_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_58 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_7_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_7_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_62 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_15_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_8_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_8_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_66 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_9_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_9_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_68 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_10_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_10_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_72 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_11_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_11_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_74 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_11_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_12_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_12_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_76 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_12_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_13_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_13_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_13_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_80 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_16_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_14_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_14_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_82 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_14_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_15_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_15_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_15_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_86 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_16_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_16_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_16_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_90 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_17_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_17_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_92 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_18_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_18_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_94 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_19_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_19_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_19_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_98 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_17_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_20_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_20_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_100 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_21_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_21_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_102 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_21_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_22_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_22_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_22_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_106 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_23_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_23_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_23_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_110 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_18_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_24_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_24_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_112 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_24_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_25_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_25_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_25_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_116 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_19_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_26_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_26_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_118 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_26_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_27_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_27_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_120 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_27_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_28_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_28_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_122 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_28_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_29_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_29_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_126 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_30_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_30_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_128 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_30_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_31_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_31_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_130 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_31_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_32_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_32_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_32_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_134 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size13_mem_20_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_33_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_33_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_136 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_33_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_34_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_34_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_138 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_34_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_35_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_35_sram_inv[0:3]));

	mux_tree_tapbuf_size12_mem mem_right_track_140 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_35_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size12_mem_36_ccff_tail),
		.mem_out(mux_tree_tapbuf_size12_36_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size12_36_sram_inv[0:3]));

	mux_tree_tapbuf_size10 mux_right_track_124 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_32_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_68_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_260_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_, chany_bottom_in[12], chany_bottom_in[39]}),
		.sram(mux_tree_tapbuf_size10_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size10_0_sram_inv[0:3]),
		.out(chanx_right_out[62]));

	mux_tree_tapbuf_size10_mem mem_right_track_124 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size12_mem_29_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size10_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size10_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size10_0_sram_inv[0:3]));

	mux_tree_tapbuf_size9 mux_right_track_144 (
		.in({right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_0_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_36_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_72_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_128_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_168_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_208_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_248_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_288_, right_top_grid_bottom_width_0_height_0_subtile_0__pin_channel_out_op_300_}),
		.sram(mux_tree_tapbuf_size9_0_sram[0:3]),
		.sram_inv(mux_tree_tapbuf_size9_0_sram_inv[0:3]),
		.out(chanx_right_out[72]));

	mux_tree_tapbuf_size9_mem mem_right_track_144 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size11_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size9_0_sram[0:3]),
		.mem_outb(mux_tree_tapbuf_size9_0_sram_inv[0:3]));

	mux_tree_tapbuf_size6 mux_bottom_track_1 (
		.in({chanx_right_in[17], chanx_right_in[36], chanx_right_in[55], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_0_sram_inv[0:2]),
		.out(chany_bottom_out[0]));

	mux_tree_tapbuf_size6 mux_bottom_track_9 (
		.in({chanx_right_in[16], chanx_right_in[35], chanx_right_in[54], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_1_sram_inv[0:2]),
		.out(chany_bottom_out[4]));

	mux_tree_tapbuf_size6 mux_bottom_track_17 (
		.in({chanx_right_in[15], chanx_right_in[34], chanx_right_in[53], chanx_right_in[72], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_2_sram_inv[0:2]),
		.out(chany_bottom_out[8]));

	mux_tree_tapbuf_size6 mux_bottom_track_25 (
		.in({chanx_right_in[14], chanx_right_in[33], chanx_right_in[52], chanx_right_in[71], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_3_sram_inv[0:2]),
		.out(chany_bottom_out[12]));

	mux_tree_tapbuf_size6 mux_bottom_track_33 (
		.in({chanx_right_in[13], chanx_right_in[32], chanx_right_in[51], chanx_right_in[70], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_4_sram_inv[0:2]),
		.out(chany_bottom_out[16]));

	mux_tree_tapbuf_size6 mux_bottom_track_41 (
		.in({chanx_right_in[12], chanx_right_in[31], chanx_right_in[50], chanx_right_in[69], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_5_sram_inv[0:2]),
		.out(chany_bottom_out[20]));

	mux_tree_tapbuf_size6 mux_bottom_track_49 (
		.in({chanx_right_in[11], chanx_right_in[30], chanx_right_in[49], chanx_right_in[68], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_6_sram_inv[0:2]),
		.out(chany_bottom_out[24]));

	mux_tree_tapbuf_size6 mux_bottom_track_65 (
		.in({chanx_right_in[9], chanx_right_in[28], chanx_right_in[47], chanx_right_in[66], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_7_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_7_sram_inv[0:2]),
		.out(chany_bottom_out[32]));

	mux_tree_tapbuf_size6 mux_bottom_track_73 (
		.in({chanx_right_in[8], chanx_right_in[27], chanx_right_in[46], chanx_right_in[65], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_8_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_8_sram_inv[0:2]),
		.out(chany_bottom_out[36]));

	mux_tree_tapbuf_size6 mux_bottom_track_105 (
		.in({chanx_right_in[4], chanx_right_in[23], chanx_right_in[42], chanx_right_in[61], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_9_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_9_sram_inv[0:2]),
		.out(chany_bottom_out[52]));

	mux_tree_tapbuf_size6 mux_bottom_track_113 (
		.in({chanx_right_in[3], chanx_right_in[22], chanx_right_in[41], chanx_right_in[60], bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size6_10_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size6_10_sram_inv[0:2]),
		.out(chany_bottom_out[56]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_1 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size9_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_0_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_9 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_1_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_17 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_2_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_25 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_3_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_33 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_4_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_41 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_5_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_49 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_5_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_6_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_65 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_7_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_7_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_73 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_7_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_8_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_8_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_105 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_9_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_9_sram_inv[0:2]));

	mux_tree_tapbuf_size6_mem mem_bottom_track_113 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_9_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.mem_out(mux_tree_tapbuf_size6_10_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size6_10_sram_inv[0:2]));

	mux_tree_tapbuf_size7 mux_bottom_track_57 (
		.in({chanx_right_in[10], chanx_right_in[29], chanx_right_in[48], chanx_right_in[67], bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_, bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size7_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size7_0_sram_inv[0:2]),
		.out(chany_bottom_out[28]));

	mux_tree_tapbuf_size7_mem mem_bottom_track_57 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_6_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size7_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size7_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size7_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5 mux_bottom_track_81 (
		.in({chanx_right_in[7], chanx_right_in[26], chanx_right_in[45], chanx_right_in[64], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_0_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_0_sram_inv[0:2]),
		.out(chany_bottom_out[40]));

	mux_tree_tapbuf_size5 mux_bottom_track_89 (
		.in({chanx_right_in[6], chanx_right_in[25], chanx_right_in[44], chanx_right_in[63], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_1_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_1_sram_inv[0:2]),
		.out(chany_bottom_out[44]));

	mux_tree_tapbuf_size5 mux_bottom_track_97 (
		.in({chanx_right_in[5], chanx_right_in[24], chanx_right_in[43], chanx_right_in[62], bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_2_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_2_sram_inv[0:2]),
		.out(chany_bottom_out[48]));

	mux_tree_tapbuf_size5 mux_bottom_track_121 (
		.in({chanx_right_in[2], chanx_right_in[21], chanx_right_in[40], chanx_right_in[59], bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_3_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_3_sram_inv[0:2]),
		.out(chany_bottom_out[60]));

	mux_tree_tapbuf_size5 mux_bottom_track_129 (
		.in({chanx_right_in[1], chanx_right_in[20], chanx_right_in[39], chanx_right_in[58], bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_4_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_4_sram_inv[0:2]),
		.out(chany_bottom_out[64]));

	mux_tree_tapbuf_size5 mux_bottom_track_137 (
		.in({chanx_right_in[0], chanx_right_in[19], chanx_right_in[38], chanx_right_in[57], bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_5_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_5_sram_inv[0:2]),
		.out(chany_bottom_out[68]));

	mux_tree_tapbuf_size5 mux_bottom_track_145 (
		.in({chanx_right_in[18], chanx_right_in[37], chanx_right_in[56], bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_1_, bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_}),
		.sram(mux_tree_tapbuf_size5_6_sram[0:2]),
		.sram_inv(mux_tree_tapbuf_size5_6_sram_inv[0:2]),
		.out(chany_bottom_out[72]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_81 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_8_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_0_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_0_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_89 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_0_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_1_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_1_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_97 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_1_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_2_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_2_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_2_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_121 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size6_mem_10_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_3_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_3_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_129 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_3_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_4_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_4_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_137 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_4_ccff_tail),
		.ccff_tail(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_5_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_5_sram_inv[0:2]));

	mux_tree_tapbuf_size5_mem mem_bottom_track_145 (
		.prog_clk(prog_clk),
		.ccff_head(mux_tree_tapbuf_size5_mem_5_ccff_tail),
		.ccff_tail(ccff_tail),
		.mem_out(mux_tree_tapbuf_size5_6_sram[0:2]),
		.mem_outb(mux_tree_tapbuf_size5_6_sram_inv[0:2]));

endmodule
// ----- END Verilog module for sb_0__1_ -----

//----- Default net type -----
`default_nettype wire



